��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��E�a� ����q��@��[��Ð�F��l��>����%ܬM �<;�#�V��CP�r�㈴�)��i����E0�|�� 6}bB����j����Y�}�8sB��Xe��N�#V8��ѯvaE\�%A J�L%	���V`z��@ND3��]���b�Z�j~i��?���$H��3~��E����;�^*
��Yg���SC���~V5H<z��83r��v�$�Z��j!����a�q�� F�;|̕�Li�����PZ\�C��sfY7e�����S��^Y�h�}7�ӷ�ۀ����6��*4�U	�u::Y��h�g��g�Y�%����H�7��h=�Bѕ[���R0�.jPsǞx�-�����N�G�QD:ڪ��N���Y�S����b���9Į�o�ik9�"� p��z�m[n|����%T��8��7��������~glF����-�G��2;̀��������5m��fT
����� ����n��'i��YAH$)G^�r��&���Q�4�3����BTv�;B�<�4�&8`C�.NzĀl|�|F�:�?���Z�c���O<z�Y3F�_�$Y���L%��گ\��7>.�^�@��� ��<��;��+0�D+D5\T _���̏��8�T�̾KIadH���m��*���u�]M6�PV!-�әc�?�A��O�pr�d+�}1%_؄Ҩ(y�A��l�_�=��+�c�X�1�f~}b��]��U�]����7��~Ǣ���е���-��{���p�3m8:���jTL~�����a+���gh�ir*`���!a��Ql��sh���`���B�=���_���ƶ��� NEU��y��#�#S���[�q�����b������D��=�uc����(tH8T1[HY,�|�1`.:�L����!h��B���B@2��.��w�
?����~�%_��$��R�
3[/�����-�y-�?|+Æ|V��F������r�;�c�[ڟ�u�1��˪sᲜ��\?�yTȲ�'8��Z5���s�*�y0i���|T���"��/��n2�}�-��l�N����,EkÝ}�q%�<�&oo��0�CQ�T+0�$�>�������k�dX8#oG������d����F��?�� �<�"��؂�o��$:�+���N��W�ƥ�kܰ�(�C�'~<���2邻T�W��>g��E����%���^�SD��fc��$�H�}�g��ٱ�8Z��ޔ�{{��*��� ����]��p�C9n�$ԛ��;5���m:��(�|���<��$�$�4���9�_�6q���Vғֻ�79��+M�c�,}��d�{M�>�i_�:�8�����s��>@��Bm��pM�E�k�	Ѫ_/[7���٬�3iu"ķ�9l�=7��"E���ׅ�z[��?����,��5��,���>]�G<G�b��ԹE��؛�v��EӃw�A�=p��nwH#}��v9�Ԧ�̉�>��z�-����(��0t��v@��#����� ��kx~��D7�v�[�i���d0O��J�(��&I	�:c$)�����p�(0��
k{'��}�T`�����z���������>���B���Qy��6�O.��ڱk"�A���ɒ���g\�*Gq��C��h����-,�VKm�����(�2}����K���,��)L.��R�T���ȱH��%�{`Z�JW�D�f�HF��4w���D�#�T7�<�+���4*�7�1`3�ueZ��f$k�-����w�P���%cѣ��N�X?u��u�gN���{�P�sc�a��������.��I�Em�@H��5�E:���:h�?���M.p��z.<��p�*a�F����r!��tә�ùux7��o����6�sp���Ը��?�%�g��.p>_�;�S���JsW8�3Hmu�2>��$M� YeU�[��^�o$l�z��#��(�e�Q�J��
���>�R���qMP��d�*u�99���n�o�����V�<�[v��_�g�/�dS^�Uќ��+��2ȃh�y�>H�F{���NtӼ��1A���o9)�W �:Nqc7n��)�Q��qJ�/���$� I�&����\,���ʖ6
4=qO��{k.k����")������D�� ���W��i���*�0����T���n)b��F���rD�q߯���:f�"}-�V�Г��b� Q�1���ա\ �����`�G/�2����T��e�Ksqm����Yz�7ʼ���Q
��x��	�@�:<�����k��'v}��؆LZX/VMn����Pd,�6�ɲ����z��h�`��w����ō�+�0`Y0��vHUS��Óf-���G{j�r���7-S^�tB	���u�"�%�'b<�W<��`N��k�L�^6�m�wK�-"!��1�~1͉�G�r�~���&/�V���6s����ap5�n�t�9w�n� �k)܏ɛ�l��@2�\'��n*4\Ȁ�\���+DT-GS�:1�7����!��~���I���I�x�r����d�.mб����A@�HF��5Fo�k*��V��dG�b�Gk����z�?� ����CX�0�����G���r����Of<֋��0���*�a�U9�l��H��	�a 3���S������"��>��v������ߞ�!�E�J<LN4�ڽ�#L-�K��C���!���;�>a��c����
-*~R
˔���������%���q?m�����"Ln+g��(o#L�G�|Y����--2�-w,��
3��y�iJN��:u���Ʋ�}������!��F��E�����Ȇ���g��
�b�A W���;�E�����l�'�[5^Vw�4\9-��f5�Q|ܼd��8�N������ :��S�1���-{�i���);�²�U_#H�d]VZ�Mm��Wa��U(р�~G�����
u�e��n�G�J�n���+IvT~Ħ;��ӷ�&�B����>C��2m�!���{��H�����ƃ�j_����~����[��d�&�K��|t>�:D4�������	��� U�#�RvFz6�����t�^��|㉌���bVo�3�W"Q-6�-��u@���m�]�cq��:��PF)|�7�.�ɯ�+���J <l^D5�>__�f���R6"�MF�/���L��8`{���>n}�شI�l`a#���J��-؇�(�a{���A��R퍠e�i�zy�(J��k^b�N��<�ٌ��N�x9�T�}þ��L�<dBi�D��{��w�e��2��֛�i4����6m����4Ƙ��|�)=	{�2�`N��
|�_�g�	�5U���"�� g��J��V�)�vqVZ�P'���K`ųY�S~����
m_����U�}>�K��L	�d>�bZ9N��<F+o�[�W1��誚�Y���K1�>�Ӿ�jHɝ�P�sc$v�u�JC[@�+����g���/�Tt 8���cE�cRį3L���F:U۸k�H�M�? �(��ő5d~笧Iw�&��!_r�o��1��ɂ��<��w �Լ��si+Ӯ�[O���-߅�y�ڴ�W���H�������x�C�q6*mp$�7�[���2��4��Dw]��e8:���|#o˭��׾�W����dIĀ+�R���f�b��9�^.*�u�D�Q}��qb�%j��S~TV}����s�SÇ�Zu)h�&?A6ֵ|Bi;��ս��'2��"���ʒo/����ɉ�Dd�
�n<�m�?�E�<NH�����!2����ΰ�������o��45�B��.~Br�~-��)����ɎV3�M�R7�f�����˽��
C;nN]F�/�}aK�nQ���C-�Чn�U�0��&��Q	��� 	x2!F���J��/�)�Iz��J����<�24k�Ok��4Uʠ���c2G#����.^�RL�Dd<��1ml�k��{+��/zA#���g���vtq�v�O�N/i�]�[*��J@r+����/T��X]+%yR7І��� ܆.-B	�嵫!�ͤ�Ms�Җ�U/��$7�M�����W���Ų��^)���ޒ>*B������ �W��+�M3'b�<��]�ԧ���v�F7;�?N��`�r>�/(���i��irQZ�!���)W�s6<�o����jd�]K{?�(=\�QQ:���2u[泋Lt��Y<��|�P5~�6��lD�L�P�`ѲE�<kUsC���g��T���2��������e��o--G2��3+�������&�>�j5VWW��8<�KBV��d`2�
�
�mn=w��\��!�!���4{��PB�?�ܨC�Pv�ƾ!����ݞ��Eš����؈���W�vS�9тKY�G�f�e�`�L�c�n�@�fu�>@��y���,L��A�TtJ>�/��^��ݴ�j�K�7�/OS�)uB��M�O�)*r�3}I�a�un�c2�V:��/�L�'��?yp� �ṁ�g�(�9�Tpf�(���w��Rv�ȝ���
���c�h��3�婋�&��uwWc�y7�\A��^N� �]�-&+j�=ь�����8�T�=U��w��3���6ȽF�X�B\q��1�Q��Q���]��RĮ�P����'0[4v\��[&n�Pnl���$Ѷ�fR�M�^��PL�ϳ������_�E�y�d3�&�z�z/V�5�lm��K\��׏A"���P �zG��/�~v$ʨ#z���Y7����R�m�5>�lIâ�eCh���ض�̗��8-��mELˏcb��=��s��A�j|ϕk�̴���:����E�Hƻ�6ʿ��(�	E�y�画�_�"��r��DBQbDP8ܒ�$k'�~K�4!�!���j�$�K��Z��詭�:����B`�\�>"HT��K ���M�a���9:����Q��	B�ދ	�x(�~A8�g��t��T� ��s َ�z��Ҿ�+\�j�]��f�1<��B�6��Z��g��0�YSTU��KE�h�[1�	���ԬoF����u��� ��pUd�hR�#��7��2 ��x����o��C��-�	��ɸ���ܦ��J��M�(ц���XJ��V�@6t?#�f6I��ay[�B��^�9Ʊ������LJî=*�f�Al�h����~
�vb�8�K?W��Nկl�\�b2��I��T#QΣT���%�=��)L�M�$�\M��|r�Ҫ�ߜ��f�0{G肦|�~�+iZ�iͿ�8���F��#�m�{y�+k�v���W.�8���q���C��3��KF���#�5/|�؏wc �]۠�*Č� �\^�+��嫖��X<Q��9�7T�2�n��( mf�ŵt^i���(La���Y��&v"�@1��3v�lE�5�R��I��#-�JaG�Y]�[�Ħ�Ӳ ���@m�xӲ{$y�m����?X��C�20��I���+x��K���b����@����;w!Q)���A
nt���T*��9�[+~)s������8�>���S�c�4���zS��ah�mu�[���*��&�J���uE��߫pg��'r�[�ڕ^��k�D
h��9�����Iϋ���vG�������2�k��Z������fG�q�
ժ�~���u �{��k[;ǻ!1zKK,K�@�f�z1��$�3�i=	0~������r?�3�����������X7���')�#��~6�����ݾ�br�L��V����J�
J�o�A1:b���ۊ�%dI�1�.���ln��C�%��-yg�I�ͷN���x�>�o�=PϹ�@uU�8)����xA�ZO'�+W�qtFi���[v]*I��ӄ����L٧��6��s���9�(����th����b6���"�ZXb�ڪk
Ȁ�\��1k��:�Aڵ0ܰ�1183��/(Q��t�SJ�-p~a�Q�$V���f�7
]��>չ,ߟ��LJcN�X1 B�>��F>�H"'�60��9�P�9��H㽳�YV�T��QX�����7�Jh	}�س�R�%��J�zJ�H����#��������
�8i_�eP<#�qO�Ô��]@$�t%��B{:�:�*W��"��{�B��D�'RR;��I<�T�	#�ӢV��k^P�������%����H��0�6��$��I�g�$�tJ�ͻ���H��=��u�kkh�|b��-��.F	�N���Ї�F"����l��E�hb�ǔUS�Ō��'��.Fk�z��O�*/����6�U�)�� 4�HV�4��3e��&��"g���V>�H(lsC���<��Z-o�{�j��+/A^I���ֶZ/)��Z���R�g���d�]��	d$����q�u8х��I�v��ZKR��8��ʂTA�[3_y7 �~�JN�^���f��Ŗ|'M�d�6NB����#�4>ð��p��	�ed�IT������}�>�~N�\Zp�>��Z������+����O�^�b���A�J$l��v����8�	��vȜ���h��s��r;L�Ѝ�:=v����L2����칪Z����R߉�!��
�~�1ԭ��^ʥ6���6[��Mjw���I����n���2�Ҷeg�Z��ӈ���'	��l�J��O�G^�`M�UdRB�<
�K�1���ɜ��4A��D,5�����/�U SJHs��B7�m��[dy�@�M#��!��Ĩ����(`j`�N��Ep�^��sP���s�{�-�[Q��N2ߓ)f|*m�Ц՟ȱ��������@�q�a�D�S���}��63gz�>
R�o���s(w��$b�����۹~c5}!��,R;��T���|�*�X{b����ѓ������D}_��R�>��K:)l��N��]m��l5B �ͬ�'�����?K�9���%�l�L����C�z��>�:��T���	�z���3�A�9	}�7�q^��fE<�9O�up�Z{x&W�߉���8%�Nd���G�KW�w!>���Y��DndBk��~���iF�Mw����J�ߌ�!�u�w�2r����H/C�l�!ԯد,��h�>� �8T������	P��}񳟚�nui�G(���:8F��װ�xo�����=�6䟲� ��#�Sx��џ�˲`*�t�[S��Liu��?0���E��7����[}����b�����n�n�k�y4�=#�-߫��g�:�~��g� ��c�X�
���=���KFQ>s��Z��m��#y���w�V�rE5h���tî����6Ml�Ae�p���A,�����,Q���^`A����f݆�G���H���c	�Odc�vsH��mGj\lx�G͉�m�#QP9�E����F2��L�#�3�@k��k�-0�#��| ��`��%��6���ծD�0_o�9�1�C9���ދ�� 	�3r��7�Dm.��ǄT�ǷF5��k>��t�����Rf�����p��Fy����V(�hb�C[<мW?M�q��+�m�����L9�4,I�XG����Ψ����z<�34�:v:˜�'�SņK�vLA(��"�9g��~#��� ���r>Ɍ~a�̦��<s)5�z�����^/^���zGƎ�{��WEm�z���%��<��i�@�G�vO����)������k�&�6�X�S+�c���F���Eo�M�͑N`"��q�ln�s�����e�FY�y'W���~��YNm�D{ў־w��lq��R���� {���������ë��ZH���+�������sxB��:�LSlԹ���pK��&�S�[a���(2�*�Ǩ&:`S_��:�ϛ�#�=�J�8=AszL\^7Z��9�m���"5&� �S�۱/+XΥ�&�WB�'��׳�0NcfѰ�i��������+�A�˂�Θ���f�u���P
�^�� �㴣'��`<_	m��rf4��m��e�P�gf_e�az�Û��L����,H�íЇ�,S���3?����&y�~����@�ˊ:�j�{�Z��;����?��ԭ�j�ݧ��{ ~�i2��˜���{�i��M����(ܻ�Og'A�����7��`�v���2Tl���x�ژ���y1��$CHu��'�,E��'a#�c|L���J���S��As-dhalJ�	3l_27��C��f���m��F��,c2�M��2�+�ș�0���`t&�1�Խ��:`E�'1F�Nk�_x�ʦ�MG�*������s����3�I�wT��A�1��q�R/s��J�{�4w�-kPM�f,��썑85��?z[�.RX7��� 1�i��s�A�MZ���ſ�P �ײ����:�)�+ÜWP��m.�g�(t�g�`։��g���W9uߡ ��0�t�bB�t%d`̵�>�{�?�b��ze�d��5�=����H�����+vd��0TZ�^����}�7u�G(�b*�~d���7�w���$�"%�����;�w%Lq^�_��p�
l��'lRj���3@W�fu�Wܓ��{X]g��׈g�
ur#V`1�w�o��_
tMeK�иA�d�7�a�zX7�0���1 ��M�&�>-E�:�C(�t�I�dft_�%�a�@,���I�r��АR��-���>'�*z�6��F�c0>Q1������W����~v�j��2�]���,�qJ�h��Ә��|(�'g6 {��_+�,dR��������j3S�L0��aG<_�!B�s�+^1L����.ۂ�%`�aK{�l&pz�r��}"���y�qZlw&��p�Z��&~��Pz�����vbh�cc�HB6�>��l
���˟s'�K(�.w"�|q41�PԼ��]k"i�Du�P�r*�<}�<ݐ�xv���o�����=�#��8���:��Ƅ���2�G؁.Ap{l���?��k/�)���z�Qq�6��Hz�SI�f�N��&»R��l�Y��,�N�A�)%�QM}��F�Dř��j�M���O3W�	h]È���� �5�����U� �ٝ5���]�[�x���'S\(�/�D2��jf*�ͤţ|��j̣=]�g\�z�#<�
j$U��?�����)�����X� ��t:��@!H�#C�;|�>5���DD�'��5��ٛ�Z��2h����Kl�M�A_<I|�}�TJ[�����e�c8i}�3=;^_p~U8s|���dܷ�a���$�.,���e��z���ҙnvj���b�>�z�y�'�A@]�c7�X��X[5:��0�92Y�wW�a���F�O��%e�)�]9�JcQ,���@:�-��/)h3yx���S�Ʒ���Mh��A���c���Nx�m}gU1��m�v�ZDSPi��
��-�	����h5�7��~AwR�̄H<�M�g�rAdm�hP����Oc:k�'B|e�9'�~�^��	�1���A�/e�����z�Lβ�����h�38���:+7�C~�pޓҰBhj�+�O��u�옥c2ϛ{�%o�bP�t9��BۘQ?3w�܉��6#�����_��J��g�Nu��[����O��y�6���b�l���*(�4�B��YW�q���]Pi*�+K29�q��^c��6�)�a��,>�ʚ�R�� �dCv"�l���$ܻz�&L���)�1�#�m��o6;���X�=�\Z��"tPN˓�6�mh՜���?�����|�ќ��M=�/���B������D���G�R
����?��A�^��%��n��&2P7_?�5���`����.�q����}?���K��]��<�5$f!|�`�l���.�$�o�j�!��b��:aAR��w"���Q��;x�H�w�z)4�;�rl�	nZg�@�²�?<Vi^�Џ��JX]057���&Uu���|r ����~0F��ϑ�%��<m����~y�;���"�y�L҅���ٻ�!��1��:�����Y�#\7j"rr�"$���۾�����޲���W���i<d&>����[�� V�u0� I��prU%Y�j��8���Ƀ�h�˨���x�5�(��m-'/��h���YdO�L����*�a���6@�9cVmUIO�\��C|a�NX����G�R ��WP�˰P���L5j�2���=`�6�a��%-ߟ��a1:7�W���gO���(�Ul:��\(��o)]�B�r�z�Υ��+���=���ﱲ�)�=���|�����7�l��j�x�"`�O����x[��w�)r7�g^l$��Po�5���sz��AtKz�3'	|�-|��)���%��w��)���>��.���xr!���d�ܜ������(�R~0�u��������a�S|�J`U8L��;\�jޔdu�wH"*��qeg��0p��$�M�*���ٚ}&����D���fb�d����f(D��u��r:���Z�V��։�Bx^�����@DE�;���^	���� �:bPZ�\Q �Q�{[���]�w���[j�@�����J�����g��k�!u��X` {OR'�M�|Y�T��҉q��m	���x�đ����F��J�iQf t�^��}M��b�G���B��z���X��R��V�#݋���LDԋQ�t��s�3��ܤ��׺3�(+� '7�/0�Mm�J���Q�a��D����$f7s6)*�^�5�4���jst�;��"�����!�� %�뗢YR��cte�5�{dbyJ���!_�,J
��Hn,��0H>�_SP�0��A\h}n���e��hS[5�Q�6�C�BdB��v�HC����8�렫�g�q�0�a	�K$k�j�_"7y�'�z�t'�uo�'�a��E�1Q���BZ�����)�a�,(��k�l"��k6��݊h�����O��R���o�Пwd{�2v� ��7�ۥ~5���h.4�9�,�\�G!L�P��(Mc�����>�["������2�T0�o���L�w=hy{smDG��_w�+;�����k�f `䫈�2�/r��T���惼	
]���K U��s�����S½�Z��y	?|b���r�P)� ���+p�{v�����`�_%���;�e���P�s5�W���F��c�uER&��V�R�{�Z2�� <�Q���.A���W�k~�6��5y�vę�:�#r%Żu)�l�=�ϔr;���u�{ʬ����g�\�J����B��������@ �1���G�12��i1IN��
��Eج�,�OC;��,Ì7ҋ� #���Ë�319�,���EiGEAbĸuQ+ �/u��7��O�C�W�oN.�\�{PJ[�g�h�aZCcK�����$�h&�ں�R.�Սe�*��+���Yl������i�<��~�����M�o�&
��e�{n%�+���X�m�]����Ep���<p��|o�l<��aN$�ME�LXJ�*BroFL���[���� �#��?e�6 �/8P�+��cK�9�3iQUa�t�@;��E��g��(S i�׮-��c� �.1tGw�?�f���&h6K�1��-�wT�5�X�D�V�XNM�k�"��D�9��o�z�#5(�3����s�ʕ��ےAa�C��L&�x����e��s��`<�ʫ	� ��L��OF��0�Z:"�*"�G-�����d����u	�X����V�*�����Yܴb8���E'��Lz��g�-j��eJ���j�#�.��/�4��
�����4�g�7]=�\��UH�NQ�ʠ6�yRhw��Sw2zK݀#��Fd�!����gcX�'���4�����_��+�o0��u�˦�M��KɫNŷ��A8��#{J���vЂ3	!��b�=5d
wQ�y�P�j���w�]~��k����γ���|@P�Bϱ��/�/'����%��B��OaD(d��5
5�A���B9�w�l�w��B:H����*�O�N�ͦ�zv��1�������=1�S�8�\��Mŉ�/���+u�n~<q��v��W�f��aN#��8�}�@��!����\sj��Q4�!��[Å�â���W��a�@445�5`��뺺;;��t��Jag3ewJ� �1O�Y�v%�=�!ꤽ���	f�8~�z��[yv������>|��֫��OU�s6�~����J�������,EQ�9Ƃ9��\@� ���UU��6[�8*�=��N�v9��r�í!]��s��x_|mO%Y�o�"�#[j$3;���_ �'
��c*�����6�c���"���sU���t�ƀP�t�d�\�j��P�J�M�	�U�W�2c��Lc8B��q5��V���������p=�䤚�E��p�LL�<�>��0*b���у��k<�Q����.�~��F�414�a�KCs �ƎE�۵�,��#I�	��b3�y���Ki��F�K��F8��I��2�s���"���S��>�X���tEc��J��*��@���V�zVܸ���2�X��L!����,�9\Aw��GT4�6�ҿ��ĮŠڔ�Ҋ8^��5)�;F=��j1>�����&��|&y��������'����'�*Ľ�J�6�MI!0�fr>�)(�C'X����u��{�(��ru	���-�7�f�
�X�,�<s�KJ!�3��|Ԗ���$��~�]���i�U,�A��(I�����0^E�(-�HK���|O���F}��o�jJ���Zw�Pؚ�|J-D��(�2�`�e��
�L5~�(DH��B�h�N�9���g���M�J��|��b�<H��f�V�5��X���.T_�2O
�!�.(��ﹺ�a��e^$z-A�)e�����u�/vn�׿?�f��x��ynn_y���]��{�R����بF�z�����K��}_����_�QM����?z%��=�i�L����B퇡��ޫȠL��i�g6�����,���m=}�u�!e~&�Ғ�I ��ȝ�*�°�rT�s}���^t��ɳ<��3�-$�eg��d]̇$��$�wn%rQ��S	�Ρ��W�R5��׍Ƃ'۷�jc?����@�b~yJ�Զ_���<i�����b�t]���o��`>��LI��j��P;&~Ї��&��d�`���(��<o� ����+ˋІ�����-˂
IN\R��1ʄK���>-���OZ�'�X�?����r�`A�7B��עӂ҆�Y�a��T����J��{-��nfQ)چS�I��gD2���#L����G�9
َ)-��7S�ӓTHA�*p�}�
e�0���\#R|��}R�z��1�VpD�E�������}1>󬅴-�^�ѳ�FQ/~�e��4��J_� ���zirϹT�T����Ӊ���V���]��@F��RQ�xmd�X��fY��W�p���#�2@V�Q��`d�5^r0"b�Z�.���$�ǃe�%8C�H��j���IL7%�6�ڐ�?��q�t��@�\� �P�j]�j�6��̕Y�Sw��u�;���/��G?�7'v��BM1�f|���Lh�|Œ�*-����8�y��Ziy��^�+.�Ȁ�q�f[g�3��.�~n4��;�rAX�\:
���9U$�!�GKlS='�}p˱�u�z���s���3h����5-�؊�u����)��x�	x ߓٝ�BD��R<�R]�rn��e����i��Kg��	Q�����㎂�9��)��Z�֒�#s�h��6k{�� �(p���t?L=��Pw��v�rA��:WY^��0��wO}��S]��3�P+����K=��+����86uC�����y)�[)�:���ɬ�9���1*��ڐ7���&�c,�͸��%]i�bMN���MBg}�L����G{�R^8w�ï;�=j��xFaG�C�i�[�^������m����
�V)y�Q���YY��񳥿"���c���X]�)��0D���|FtƜ��-Q��a՛��GI��lO������l<v��@7�_�<���un��ȧa�|��2L�#�3M�D�Q6\'L��6���baj�r��U�;u�r:����/)r~R|`��x�#
�V>�w*�ء;&_�?%;`�wY����B�͵�F�oN%�#�X��p���yf�$;h�]5n���̌%(���P�R���M�=��\]e�O9-:&� �]�"�a�	���y�ߴ�cD�X
��Hm���␋}S�e(΀ Q��Q����X�����k��΃7�B�i1!F嬽�T���G'#Po��ġ��tXb ��X���G'E4k���q��̼}��gyg
�2����\igŐ˵��W�oH!b�X}�G�z��X)��&./���ƙ�/�_C��[�#�=����E-�W}�Wp7}>�u{_�xN`8'�-bgµ����8��x��l	�����z��X���lzm��8j�lc��`Z%U�A~n���ƺ��^��a�&x��w��W�F�70jA.~����}_���'<�����h9�~Bi�Mi3^�]�Tp��xB8�
�x�@5�q2g-�`��Q�D�ҥ�խJ��M&����ata>��o�)�!�7M�<���-�������χ������c�Ef-����I������h�z�@�U����y����.�g�~Y�a�YE�����2�i-�p�=^Ĉb�Zv�fN��������M�wj�����cJb��j����>ض2F��Z�&�J�l|m3��g{i���b��kO8n��d��"�'�����l�Izq�����	� \.�5^[�$ν���N����P�*�B�� E��*���LF��<���r����{m*`�4挲�F����8�����AyT����H��ԟ�����́˻+�[z��#�9���r��0a�ձW�z��
_�X�P?�_}-��`�2��Ո;�;��I(>8��~��O/���t4���
+ؼ��@�F�5��~�ɦJ7�OƊG���6�s�ʌʂ��*�q��tUD�y��pI���IY-I�謕���tx��+�����sZ�L&��L��:'xY>R����p>sҡ�'�Q���MxFD�ιx?�4Rμb�E��%�
�ʤ~��̴���\��It�*�&J�	޽�)��B�N�v�����
r�l<����ǽ\�V���z8����"�ih�M���LN	����M	u=�,Q��r�Gǡ[��ƚ���P_��e��cG�B%�CR-s�_ Loh���0-W�H�<ڠ2��-���?��IL��Q�UR/��U�-�+�"����Χ��0�֙�V����=�@I�D�v��d����n������P��}�u)�@��fޙ��84]�L�$Re��<����@^/�������X(���Ӽ?b����Y��8UK̚��zv�H?*w�Z�7�pGܘ�l{7FT}^y������Lp�vut9$~�A$[�fBp�g����iD�}��t�C�m�1���|���V�;|���}��c:�Y����OV��j��t�0����>>s�in7&��
���u4�I�����A��.x�+>3c$��Tz������r@�6۾�s�"���$+u����Fk�Y��=6o�Z�M߉4�h(`��u�f��|�4���3�ؿ4A2��q��<n=Ot`��P
��@\�借�L�65�'�]��Px5Ve��keA���7�T���.TA�~uh�^����͙Qi�aw�G�gYQ�u���@��8�T�]�lH1వ$��_�`D�R�υ���Q�Z 4����7���GI`����$�G3�E�I�[_��N�ِAO6����_�<&?����ö���Mծ0N"6F��8��K 9,0s�,��R�,(õ͸�	,׌��R�Ù�	,�~�x�]q �_`��-~SѿoK"�b���
��Ķ#�+��Ttb���%.�%H��3t�����Q�U��(�+�,�xws^s%U���P�!o���/�1F�Xp�j�/
i�F�u��VM�p�w��׽n��)��޹磺*�Sɱ����+"@
�7%�u[����k�(E�Y^.�)�ׯ�W�!�o�FK�l��b
n�O�ɢ4C�b��O8P}��)�咟0c�ީ�G�Z`���*bD���n�B�z�c&{�Ƙ����Dǁ9yM6������T�~�;.b�w���������m欜�{��>�Ǥ��c���[1���:��Bs�=�i�ђ�w]d���}�)��L.؞jRZIp�%�k�Z�Ns��~^��������a��R�\c���SE�bLBd:mm��R4�)v�6�A�"l*�i4�(��_�&��=o��Yufc�ɴ� ���9�����n=R����~C�g����L���WA�1��䢺�2;O(�ܖ����3���Ɓu��Z�7�R\Bɿ��0ci;$V�NK�=��R*�*�c��<��A�*�>Br%[�6�_^$�4�
�Ӆ�r籧=��o�vS8���~�,�M��B�{��V�v�3�� ��e�M6Õ$ͨ��hNd��1N��9]��]%X)�V�L��-x�ي�pO�1�f>Ɇ{�	:l8I~ղ@�Kx����~�r�yPW/���9�2�½k�`|���u*#�<�Ҁ<ޟ#�us�P!�N���a�d0��qR�)˴U_$��T��CMV��Ԥ��dQ�յ&H��]��(����QU�7B�e�T@��!���l�Vb(%U�19C;�w�?J}by�u��b^��ɵ�]jZGmzMv=b��-��Re�(,�?z P�Q��o�����1)��6��B��Q�tg��W5�e��������Cft�P1ڠNa�����C�W�#�͑0v:t����]�[���ˠc�cBn��|��J��ڜ�n�JFV��6q��A��i���^����n�2�(�Q���'����[�8͸j~�+_{����+e� �A���ˡ�Ox��;Y�������ٗ�H�>��`I��y@Ͷ��t
-
2h^�آ���ns_)�	�$��ɚ�n�������\A�)�<���$1ԋ�}N%���S[FS��C�r�PC�m�ejM/�9����B�'���WT6��ꆀ���y��k�:���O�m��z�� �\[��`�P����<	��fd˒��hɎ�͚�K��������B¦ZM��W�d���n��ZSn-{����������;�ajM ����юb���"��=�*�y�P�����9�:MPbQ%��e�7�h�^g��0������|��&���ҹw�U�����z�ñ��h����<�Y씡��:#��z��{ ����� ���md�ONO���)ґ��?���٧����<��?���T! ��2K�P�o%�C$�_h��6@p]6b���pX^Bd���c���@9.�%�+Xt����"D9�P��F!w����>J�}�M�`�l�0+��v�f+�u�i�=�w ���U��13ͧ��P�L>�������Z�Z��ur�*�r�/A��hC�o��%�݀$���b�gw�D���$io���Y�nCu-�P�2��F�\.���թ^���N���<�������
�:��W���c�����s'Б4�mD�� �y�0C��p0a��f�G�|
��Kq���n�ڐH3|}U�{+��ۡ�������I-���mWu�|�2��8�9��dh���K�'(覨sT<�4������ |!<qoE�4E.F	�YE	C�<2V�q�M3��a��n�P;�C�l�gj�t]�R �J�?����;f���-�߻��6c.�spt,���3w�R��K�ů��X�������-\@
]�޼�AU����f��T���P���m����A�#m�(�kw@�I�,U��n�� �ts���A���5���>?����h�Ot|6d����չ���ɧ͙������#L�'��KFNV�����k	fK�X��FO�T��Zi��}A�__�'��Q�;���(b�J+Q#�BK�Zy����G�V>��Լ �F���`���׺��w��C+�t��R�"8�4HQ�)�ٞ�qу5�^hy�oNt�Q)�%��65,�O�|i���y�Ԧq�ɻ%�k��*��������	S'����H��`�;�
re�;�q|�~�y�zz{���܇��_��"� kah'�e��V�০@%~�P@I04�u���9��e� ����m�m�����=��P�(�p� �Km,�j^k FK^"�@d�NW�+��y�Y&�n�f��I�?�;��f4U1pJn)~y+C΃'@[���S'�k5O�c�%u�q��Ğ�ͷ������S�n�ݑ#�&�
�+�ǃ��A�1�$���ظ-K]���tX�C��9��A���ߣ3��Jd�N����խ��e<�\�}����"���s"�U�����9����Q`]X`�#X��Ǹߍ{���A�-\Rxlp ĻPU�_I$��(ֆ	M|46�>{�a4 	�K�
HW�.s*��4|I����>���BД��dz�K��_j,u�[�fL��h�kZ�$83"����S���k���L��b����Dݨ��og�,g�T]��2�r�:̌�qfu��o'=V�pk�x/�qCf���0#!_7J�Jv��Q�o�-�5�&�M~���:C헸¶*���evK�i�����4M-1�DxQ�p�fQ`�yO�N����f+�nhZ��e��R�37�>����\`#���SwbR�/.�!��[�l����(;6��=�n�	9A������i�3�z[�>u8�\�sM� ]���W������ֆ�Z��k[��7�r��7�"�c;.�� /='�◑@6]e�����<�Hj�4F�}2�_����%�@W-7B�+/jq���*�n�nh]�E91K���<���T%�}w���U�Z����P�	Ǟ�m~����Ӫ%�ԡ�� �;��e��f5��P.�HǏ��Z&N]O�=5V*k�a�c��?��v�(���o'x��o���O���o��(Ӹ�ķ�_�<*j�D��nH4������[{Q'&>x�U�2Wݝ���L�;/v[�� 8Mf�<���}��1�מUY�F�
����)ä�ݬ�絖5�M�Txč~g���t��Ր�z�M�(�?5�"w�M�tj"ԝP��E�5��v����w���]�����1�$<�ކ�h.�M�9[�y�[���U�"?���qګоa*Q�;�h�\6����kL>_�O��͙N�٫$��dAs�̎�l�f5G�p�H�� �")�+:[�n�����r\F�b,�f"�ÿP,�}����V��Q�X�	.7s˭(xr���1=�?��~n5��ʞ�TZ�}�f���r(�@�!#A�����&���k�S�zÆ�'u!�e+�I�B�S�䲞߳��y�QA+��:�K��̽U�A3G��/z���f'��SJ�J&j���xl-BN��{�`{��L��	��tcu�/��2p>}((�m�S�i�mLѭ��-���Y���)������+�;�p���T���<�L 	{�� 8�G�(qN��j�����՗".���SW���\P��5�/��˛0w{�1{� �x��]g[��v���[�vr��^�Rm��v�߷�6/w�5Q�u���'&�Rs,��o̺j�ilV�~]и�_�*�u�OqY�?���)�,�����оc���;�M;�L��-m���a�迬�s�%�Cnaa[[*nD��"��8��l�0�*-�}�i�?���LMH�QR%d���q��?�k���M�ř�b�=U"��ȬM�Ky�hM8͗DAt3��wr�����kH� na�2`�W ���¤0�'w�,�lI�$T�r��LU�5e_Z}�_%��x�j��ͼ0���5��_�)3���~���J�����5����"Z������槳^0����S�H(xŃ����1�"����}0A!೅
F /���z��)of���/�~p��,�֜��)��<�iC�ҷ��ӯ�Z�ა^��z��1�K^�_l&dw�E�rLuY�~�R�|�7c���Qi4z�qa}����q�@CЍbB�F�/��@�e{�_�#ҒC���g�;T�� �'�3��P�!��\�7@�'��
����h��I&n���{��,���֓����c9����]P�}���β��}�J"7�\)�gY6~��e�3X��\+��v[br��o��PU��_)�7h%�R+u?��� ��`͌:0�ۈ��q��{8]��֔��pN�ve�5���k4e�7	i:�
8~�5���y�3P����[DvCy�C���Cޡ2�j�āI(c�\�O��D�ԝUO�O�F�	�`���ʢ�s@���S4;�^�, w@��|-z��`��� ƿ�+�G�8����h:=d<�ˉ��O@6�l�b/�D�.D<#��X�Y��If�C`�K�fK���aA�@H�a�Y+�Ҭ���t��ig0}����o���Lq��.eߞ����F��tro�:�!�N�"�n��O�c_��惙�ʘ��*Y�Y)�$*@"����G�Di��x��"��� bA�#!> ����y��;2qo��
��4 ���J�?}�	;�4��$ʻ��Lc��
N �F�t���}񚧼�'c�4��v/�.�?� �B=��y�t���rXI���(��2'fD1Y�E�9�=k4)Ǣ)�<Ԥ㊱����XE)�׀ӟ:htYd.)	1���L��Cqv�-�r
�ߣH����_68g��-n#k�;؟�Z�'�Z=�O�"��J���D�`�W�T\@�����k��3�.y�%�+��,ꜣ�Aq�Y����xpn�q�:UV�d��$ۍ��3�yѦ��n������G��|�r�6��wi���Ŀ]����o��!�~�=��_��X8��d�)W�c�\������z�Y�.��e��?Mp i �c	����3���x�깓W�n�^O�~_B+�/4ƒa߁��Q�#4�
�iyҔS�2N�n�_�Y|ȴ�s7�jmV�O�b̶O�\��Lx��'3����:�@����K�%A;������3��=C���$�mA�}fC/�x4v�w���7wpY2Q;�G�Y]0��Z1�̉-��>��?x����HX�w�0�@���iq�V�rPb 2(���
:.��*�����q���������~k�|��B�9ߛ�j��h��ɿ�ʾ�r#�=�:�1F
<��|�J�Plj�KSa�+qїGkǼ�7��y�+����u�?�P�~��E�ǜ�Z<>��  NN��'l�P�(g��Kf����q���tM�d=�N~M�R[�Q� ��tB^k\�C�z
Z�Ƿ�pj�x{�@=�Np%��K=�ȸ��A�S�؈�"1&��{��vřk}'��L��'/�aN0�L�:i���-r���C ���)P+��?�'P�!�� ���D�����fMH��f7���q���'b
�.�Abt�%�KAS�;2���|���wJ�Sl�H]����{��&o��3W�K���K/���ћ*8fk0%���:P��M,0�v5���9�B��1&���%Ȕ}�M����f��3���xD/	)��I[T��OG=�6;�*%��J��ȶ9	G�f��Cܹ���Q�wiVJ�՗]ȇ/��!hnR�1��AeE#2�F�# b]bW/�N�l	I�$Nw����pK\���(�6��i�������Y2�Q^��� �ԎU����r��'�UN�t 6��ƅ�)+t��Zi�%��(��r�c���!�Oɬc��3fUh�	����5��)�y4y�h����U��GY.SƱe����:����>��=NM����!_�Z0�Co� �]���*�e�D/�	� �yO��FJ�-&��'�$Rڱ=�M�]nu' dpKu�AT�9^ ���;_� ��7H��SD����� e�H-2U"�3�W*�֝���n&̭`���m2��X=<�Q�2�֙c.�n��N ^�=��B���O�� B��v>3V8�#�&j�]�W]Y7�\�"�4�9�޴t<2t�|�~�5�)I
��&�P������'��BT�U�4��-�.ũ��Ҽ2�üe�Ih�0Ҧ+ݢj1G+õf�5�W�M��7��r|���ϝ
��C�2�O5����v]�l�]���^��c,#��q�Qtü#�t6�Yu��0v84���"P��)M6�O��Ǣ.�8��둿S����LH֋������8W��u�,w��X#rvҗ�4�t�& ����Ǘ�|lu(��g�Fo�L2�=�W_�!h�����f58���n�>�Y;w�i6Ɩi�w��}d��H[�2��6�� �ԩ�2�&&�vD�Z�]�$��rP�ܒ����Y�E�dw��J�Y0�˻b})����B��i�ڙ�:��P}�W*�5� c��ҟ��~*2.U�]bǚ�߱�ԫ��*�*��!��[j/֒��o�{S6�Ĩ�>��g��F2n�A����{�����˶��]/<]ؕr�Zk��<��{���B�YT�Y��G���&�^7x{�~�<>Z��s5�	�`����6�QWX�Ŕ������eR?UF
3('Q�dj/�DdL�*�Z��@pL�C�}5����{�a���C~�6;N[��Oc�I{�g�K�i��a#�zp֟Wp�t<�.\i)�_%A��3�� )�2Ͽ�Mڔġ�� +=�@~;��-��t���V�'@;��M92JN	5����T���	�w<�̂8s{���kZ&��%�� h� ��^Eф�ͪ��C)iRm�>=���S0Нt$
%;ժ�\����@�ߨ�3@���`=Hw?*)��Hףr�>z!�%< ����C" =�?:�x�m�����~��4E�l@�~�h�|�Ti��p��MC~͕�d���KG0�#_Q��U^P��0�Ku��y�U �<�����*å����u�.�T"@�� ���E.���a	N��5�^ l�ї���Tb.�cc,E���/k��o~�bk�1EpX��0�� Sͨ��jp��
Wّ��w�p��'��s-7��7|o?<J%�G)�SKu��y&�[�x�O&mэ��f?h�쎚;���cP9�{R��58O�.4�_����*�]'�T��l{|/�qȻ|��o��<D��MN�Z��e3|��,��$MZ���q��+������Q�f �;X��h�6�?<��E���&�)W�68��H����({��%�k-׵� ����(�����K<a_Ř��"�ۺ{�B^��w,�,��k���Z��%"vT�ȅ������6ڠ�����ǁT�]��0����KͽXc@d�5s�u�L<f��o��w�E�5�'� -��	�I�����N��i��:=j�@2�Ji"C!2e0��o�&s@\���l�aO�<�N͔���6a ͥ�:^�HW���WO�gS(���E��XάA��r�3!:���7ý���!�[J���{��	Ɣ�zNG�����x�go���!%ٺ��NGv]H1�!����E��8%
�"��0퓪�#��|�W[2������;ѵ�`�ϫR�_�  ��J�W/'3$�~H���_j�zCm�:Ob�dH����]�zW0�N��&Q���4�/��eݖ�G�8�	�jd��KL\��F&ʗJ(�����&��1�P<C	
"������y�8�U^�56ؑ��1���������k����'$����A�&kd��>2,x�_���/$��;B��N����2��\�J���՞�ʔ"q��Ƶ:�=]q�zA���>D��a�6�T�E[C�$��Q۰uq��q�M �U@O,�NH���(�����|:��6���N9VG�#����Ѥ� h�-�t!b\����z }��<���OvZO�����>���û/����?�E���0�o�-qS��.� >�T^ҡ�;�"3��tݱy.&N��ΎO�nc�����!��1zo�\}���m#���C� U�\�g�$��< g���b�a٩?0`�f�ͽ�.FUN�jsܒР�N���X��ҫ�a׃_t@�y���4�<�̆��X�Ȍ/ ,]�p�i
.�Lґ���/�h��!�fW���6�Fp�����[r>���:�0� �\����p��5���;i���`�	��w�L���q�!����tx�zU@f��u�1���(�hDC/1�/\���pbǤ��ʩ��}�~d:����<���I��D�PWeȁۼh���o���v�a$�Uf�gI�zO��ח���*D)�y�Z��R�<�u�du�"L3�\f��z�k�8ݚ�UL���&�t����z^'��g�O�����OpS���B�]/�#.(�H���ܾ��j&��: %��S����5u-b���hKw �I��c4 �ZUz�:�]�B�l!���T��Ч��P��<�Ew��"��w�f'=�d�~�A�grd�&dKC�e����Lo���� �+�؊��ASSXboR`#�.S6D��ow!�8_�8FAu(ㅲd��G����������@������&m���j�0�0$_uac -e�o�@"���a�iKg���5ڲV�����[�<�OL�t�9}��E+-F94I!�j�
)XD����~9*oMFnd��FmF7)�$����	T�	c�;�kӷl�$��"Ӄ��߀X���Wj]�[N�\�B&ۅ��]ƭ��(�ty�#⛒�g{���{��鳈�3.d�)�ꢔ���#g�H_����8B�@D��@�>u�Dɩ�u�ViN�9W��,/��-�7�����<�i;uH���_䍾��E3K'pi�p	��r7�&���H&#ri7��v&�i/����p�ҭ�"HkQ�?@փ,�+=|�V7�� �Xns��<�{	ώn�Bz6��m����{!ޔ�r��0n��A����|��Au3"ɛ�k>9�1b��A'�cf���c�[�&�����/����)�=��r
�"���	�a�$�{ׄ�4W?�u�U�k� i8M�
3�;!��B.v8��������SݕHp�Sx%c��|2M���@��J]N�g6��@ �SP��w�H@>QHjWo�3˦V��)����ެ��
-��p6k��e"`��4�th�p�n}�Z3bl���������T5t?�!i?"hP"��F�A���e������fڊ^���`wu�R��o��f�*_
9/D�#[�5���c�/*��y���H2�H�pT#!�X����d�$Yf����ג爯��dvI��$�߇)^�0f_χ|�
<㗤�V�b�+,z��Kۇf��p9��דp��\��M�媐L�N0�rx������%�;�]�I�|ޥ�`r��N'�r\"<���:�������i��\�ɺ$Z�
��}qT��e/Cd�+ �`������9��w{婍��m�D��fO�;g��nm�}�iV'��IW�O1Ns��˻�[Q;����[�jXFD���
d�ÌD*���M�t�K삺��+��(0%w����#�����<
�Ϧ(>�s�s_c�M�i��~�e�����Q0�({���bO���wqr�]��p+=��?2�P��w�P-�l �� q3�;�sZ*��b6*���o�����]�+����.y]�P�6� ��S���s��LF���{ų%�-]柪����\}�>��ls�Pǿ6�'����Ъ�hd)���}k�7yz�����qB�A�����5����,�wJ�W���JNJn��5�XuK���z�-k��mꍋ�|�������7�������Z��w$������g�`$�g"�9=��0Ol
;d�+�0�qe6�GD��4�f	��Y,����5\"�<s��j�����bľQty��O�|�.�#M���n��ͯ09kG���RjDF��Z�+����V���=#2��tM9� �9|���3�9A�� ���:wI�{�mc4��=�!�W�'�d��J��nZ�p^���Z�\w=��]�7$挕���o.#�y\�ܺ�u��ᒕ��Ȏ0���c��v����z��,��5�b�w�bc������a}���c�,���5����q����h,yH�&��������$�I�z̻�]T-�Ҧ��'��p�<&=����ɣ�\�)"���5̪�9��3�ji1�����B(��[�E��A��b"]��.14����RV��+��vGF��W�T�z�����j���g��'�-��gf��~ ����j�l$�qC�)�2aDQ�.$]��l��f�m�-U��VA���!k�ó�W�g�P6l�i�y�J^0fH.=O�S�M.)�i���.d!Ak�8fzl�+�����}���'f��hf˴��4Q[��z�u^�����FEn�>��	�-L��閒r���[o~�(��q<&��9�v��k������ء�4g2�ͪM�f��=4m�Z8�����K��I�0�S�!p8 $�9�����S��ЪӴ�a��f�������8J�M�\�|�rZD�;�N۽Ί/X�C�����U�%�Yq���opa��ds��ahk��N_��=%k���<�2<��(}[��*��^�_7F�y|p 2���
��s��L���Cr1�ke+�J"i��Zx���}"��}Q"F��mMT�D9 .~�R��u�L��6�G�����ߴ!���^�� )K���*�O�?�4
���_K��<u��r��;UUL���.u_ ���X8b��ڂ	����g����f��V_��*��i*�`��L�H��ݥT.3g��E�H�p��+E��f���9 �%]M�SZ���5T��z�'���[F0�#'�}q]��W	�m���RXX�����MJ�#I ���s�Q5�	��p�K��Ȫ�vyK �e�w�_��,�#R�UӅ�|u�������R��^�i�T��7{{ReϢ��PU�g;P��i�l	M1���+�R���a�����	+5R���yAL	���z��c����j����BE�t���}��e:5O�Х�V��QR�Oͬ�d?�1bcs�|a)���=��x�}/�>5$�u�o3B�&�,��]�5��e��ɅTV�����욬w��Yɵy�����c�kL7~P<�SW��M����b Fy�����vkZ����H#z}ֺ)�� hy�)��:�
bVM�_N]mǌ*,��>���sq��;��aw���l�aս�7Q�W䅒I۾�A c2׮%�DCW��Q=_�p��m���%�M�Ba@=R��S�w��	L�f�Ko��4�ae3
�vT��re
�:�Z�-��iQ&_e�^?�ED�!6�*���zP�&����&���h�H�L�O�? K4a��&�M\6�s*����ic���� B��w�?*�}�f�X�eM���%�F��_�%M��9�g/��b�egA�Dl<挱���<��rG��l���<2�)��=����a��q��
��_.<|>�D�G7�������Q���޲�!��}ٯk��$E��ƣE�}D���@q%ܻsiGK����/�k�T4{)��z�]EF6/�tnJ�q�&i���IKi�c]�3�l���u�xLϽ�ܾO�~Qr�g�⋕�½fL�QK��^y�,�O�Q�C&�R�&���y/6^f��ɲA��"`N��Pq�H1h9!{��ǳ� ^r��'�	��+����)�~톣	�Ӻ@����@+E��V�'I��Ⱥ���+��vb��=S���R�x~���)!G�ʖ��W�TD"N���{4���+�坥�J��͘4���� �}�B�R�ʜoP�Ȅh�ȯ���5�G=�E�[}���������VM���l��u��U��b��f��		���gՆd��}]2;�G�(-0}X�7@�<żLГ��cL�aF(����'���kA���MY�:�ȁ����/7���rSWMJir�s����Xߦ �J���n5�*{Y��#��=��V .����;���93�V͡n���&t*��y][�g�kT�,f�̹4�`��ފ۸ݨ�L�����̭pvp�/��&;̄�t����@�e+$"U ��gl��TQA�ψ�E��e�0i0'���������>����b̃R[�xz�{	ca^�y�A��`R��c<4����,�r�OR����0�Q���?(�]S�Xu�~���q���&��/���b'B(s����a�q�N��c��:�!1fp l���m���t$�"k$Ԃ���LHuQ��ڈ'��?�3�L>�L"��~U�0�{cJ%g��ma���p��=.1��.%,>X��@�Uo��U�	 X�KB��ҷ���xQY+�6�l�n�\3�?A��W�$�����g�&�|���G*Ec�1a|2Ɍܤ����(z<��'�Y{�)��O�8+6!RǍ��11�'�:��>���E�I[���| �`��1���Ka,4���+V,詈�3eK/a��������Z�9�uR"M�@9(����dn�'z�S�z����+�r-,3��W掛0����r�ܓ�5�-dv6�"|q�0t�<�����?6~��d9��P����V4]˖�q�ڼ�يE�W���H���X�������]��3��<WPޖم��(�na��,1����c��ky���\�< >�0U-�s8J��2C+5 li�k�1��Y/��������bCW���4�1�G}]וu����7H�za=�@�FM�Qe�{@�xz����r�C���*b
Hh�A2	MkY�	md�|Cb�$�q�ϒ���#����h��־5u��n�tp)�����D[���گuAM�+�&�(+h��0IR�{��U\,Y(�)�,�6���w~��Bo=6"J~%?�!,Na�E���E?Vν��Z*�L�!t�|��\�FiWE�Y���gq��?%�*7�'�;pF(�>�K�cţ@G�<�����I�{���^q�C���=8C}\c�@��9�O}>�;(U�(���W��Ȣ5J����W^���Wܩj�E����A�d����3��$73{V�`����a �kW$N�\0X	y�@}��.�5�)�׊������������ϖ#Ǧ��XΰE/�'K�w�BT((�^i]�_Y:Qz��,��շ���lDs��}y�澐ڨ������Vg;�����i�"p���㫵��GA��TQ�˃K^�d&�07uc��bxW�Д�}lN3�K��^ѢD��Z#�γ	�>b�����5��B\4l<)ϹP�MHJv�4�<<(E�ܖq��n��̣@]_#R?U�*�wB���F�K��1o�z�͙nmF����8X�M!����Aq�fӓ�|³���"�[Ze=F3�(4���MNܼ������oBl�)K7�	R<����Ȼ\}^�]������=�c%�:c
�!�8��qiB���`�=�k@3�e�n���XAM��m2�bL���D:r^�Xz4�3F��k�~�ںTyD��'��o�?ܑ�] ��E,�����ո�}�QE�?o�f��/D���s�����
�W�&���"[��&C���S�eT�a�`<�iƟ�W��D;xF�|��󶴲O�U�=a�- QŜҀ㑓^Hx�L����5�E4*Cϫz��]���U���7�<�&3�p��L�<8�A�u�67���=��4c�{�F7�r�cL����Y_�I������I.�3dv�9S9�a�)<���۔�W[�9zI���lF7�Ξ�p���2���x���,(���C"|S���'�����*k���o�Aی���f�l����$�1S�� �� 6�'�=��n�}Mg�����b{�0��6L���1�☧��i�{�~0��a���������P^[9�=*e�}�v�0�F�Za���p�Ѽ!�P���Z<��*�n^����+���˩��z��>iW�G��'C�7%�qx]nJ�� �2B�������J��������@��z?PV��J4C�ET�xb��$j&�V��9���m2�����
 ����*t�G@���1�؇e4F��$c03�ngK#�^2����tAB��p��k�V�9�m�1���3����,Q��_��Rƌ�Ӏ�=�����벻�����#���P�=D�L'&Yn��%�H��y
y%�͡��2n���T�y��Y#������B�����nG~�N�7���v�T����^W������˙GE�|����{�m��+�a���� Sm�{ �/�x��y�O����Ɲ�QUcH׉��k��Z�A|�R?���ck�p)Ũ���<���Η�y)���l͸�������6!�7�WSl[(�6�D��ڎk&Ε\�%t�AOA��%3�.
O�>R�.��q����jϺ�#m�f�Jz�f�f8jr�,�`�Ӗ���7	�S[�[У��n�9u�}��'����yK��Ҋ+��2��W�,L��w�}�L���
lg`�����K��%�HN��z�ȳ	�R@
,p�>��� 0v����x����O��b �|�#R����� 8�^qiϻ�vT���|�R ��.-� ,v��@�â|f���w�N�@G�4Q�c����}.s.z_��JN&^?����Q���&lH�XSî]���%j�逺�ծ�ps?]����,�� ��@'ܟ���=D���m+�a��N�ۆ�vdK�}�b{C��{P��x�5z�����6��s|�X�u�{���6�}�b3�L�HM�r֮��]�:gG~�3p2l�0 ����u���A?!�T"L���tҵ�_>��_'�o��.糏�JF��(?�� ,jY��
����.�XPݍp��/���1r]M	�A�5b�J����xI�Y'	[^P#�!>ChC]�P�0�I(l�r9f���/��\+TR�>m��(�+������ ��@Ì���P)���o���Q���	1���Ž:Oa ҎŇ�U���J/O��:أ�|&��=}����?JSI�������%�K��"�����B� uݝ�f`�\[wU��l��o��[e��H�i�H� ���3���������^���w_,`B���o��'z}��阕���!�UGżv�w�[���K>F�T�AG��#3��Hd6��pڮ3�H��wEMX��E ����$��YrB=B=�����WjD�Z�yl@C����8�,��=^� N��<Y�P�-#5���n�ថ�3Y_��}���-|�����b��3Dw>f1«����;�:�$W1ݺ�t��qf���yVg.}��)�Pz�_fh��O��,<(��ܽ�"�Ax���X�z���p�&�H"c��V�==���8���l���n�!�l,��.|O+I��=9�E����I�� 3h �v�4k�m�<=�趠�t5�g�I����Z���@R	�b�RSjX<��V��YQ�A��O���c747��"�U����؜�?�?=2�H7�"�6|2@�z!�94�E������W���2�B�Xf�A�fyb�x��Gߏ�t�Xxe�#�wK�g8z��e8���K�K)_��Y����8T����ݠd�6V�(J�酻F<m���:����W!�f����7��:t� 5��O+�\*:i��*�w�g� �㬱��l�Dz׬K�u�%�z`��G��x�O�C���,�g|�Mo)"v⯷4~�Ċ��C?ĿT�$D���j�8DF�o�8G�V4������3�B�c���{E(�-*U�I;NO2�I�r���k;=E[iT�ӄK$"��j�
m	|�u�Y�b�-u������o����J�S!����ua谍�⯖�*�!A'���>8Z,
Xۺp�]t��;2��(}w�h ���W��3��,��� s�������^Sf�_EB��G[R�ԝ+N�	rҍn�r����^�4��f�QA�,��B�"�1��ԊBT^0ǥ����]�K .F3bӢh����S�'�з�C#���g�!$�!�(7e꽴ŚD�&�N����	�\�篒%�7sZh��|��0��[��F�G�?�v|�/��L�<u#�Z�[�,0VO.j
�x��$`aT�c�����8���7� ���[��Q`;x�}`���ܭZ�����<�jzD]���^�_��T��7x4��p�~�ko	��9�8�#ۤ����,"�����?4���,�{�$���1�(��,�K�.���K}��H*0�v?ą0��b3Bh�h�K��vI�6Ou=}1�4ɶ��-]��s����fѼ�ݘ�;��������7�̽7����]��|�a�h��E����_�+5K��4J���ى�O�ۊ!����r�v�:�7=���hҸ>�<�K�ZiΉJW�f>�c���؅���Y�8r�l��l~��3�4�3�+���|x�F�Qi�:D�'��y��*h�X�nP�ь�J��B�A�-mW@��YE�f}��C�e�����P�*��bv
�����݉��CTٽ�?a�/u��b�=�z�$���VW#��\A1�Y��[9![�]� ��,�P�����U�)+C/(���\�q�qg�w����sI��Y�Tbà�鵔 +@hb3W'��(ξ��aE<�7���Hj���
@j����(�9En:e�4����@�m�_+�L�rJl�r�XL�mYkp)�����)`0���#�'��fS��Q�ݙ^[���,�#��>l	o��l#Z1]0��<J��[�*�
��iIo��^~T4y������V���� ebt��Ƴ,�a��ns��k?��η�p�}bSX�-��'�i�׹4�M��o_}�i�s�r����w��T�kM�+��A(�C�Вl @І.�3O��O�ƽ�c�I�03/��"�(G�nt�!XOٳw��y�ԛ'?�����F�{�lڰҦ�_Q�Mcc����)�$�v������[X��NO�	�f@��/üӢ.�sS�(�lb[���l�������\Eߐ�)) $ "V�9�95S^��9]^Nrh~��*a%�X�� "�����_�i-�1�г���U���A=LW���RfA'�u��*#X�B����Tv�}Jr']rĶt�:&��`�iշ�6	����=)[���J�����⎒qg��"�Ɏ���-����?�_���$�N
v�"q�,wJ�0:��P�\�/¸/O��0�f;�2��ґK�!��-�PS�
A���z-;i6���!�w�[��7�`��̺C󨫍�`v�P��ޅrBY������F`{��v��v1/��T,4E��}���>/�xl�E{ͧ�~��j׎S�N���Y6dC�I$�w)�
�J� ��x"My��?M��Y'�F��?��	�q��mAZQq���Q���S�׿�|ɘ���m�����Wи:�B@���ƔB߅~��EG*�:��ꗽ�0	^��ۡ�ۇ;��~ҋ��\�[�n8}'�%�#�y���̰��Pk�Q
�3��dՃx�fEd�V�0�sI՘��/�2�"O��v&����~�\K� U�Hh�*2�gRd�+��u��[OJ�M�O
2)[;�q��|�g��$��`&Z�2d���B6ξ����R�&�̀O_����D."���(���?��l����qB��y��01��3fR����(ǖ�������~�8�"j�6��&��*|�S��ccZ逜[��:]$�0��1�d�n����LLd}:�O+�=�)��ݠ/[���sf��������_��	��X8Ci�� ������H�x�L���o�2�+��hn�J��'|��,�
���r�82;����:r���l�ZA�E�b/W{�GRM/��覹e��u �
�y���-��|��q�K�dT��0$x�������Od+���;I!	���A,�D�Z��U
H��q���g)<�T<Ke�Ϋ!�}���L�?��|�X���
GK�e�{`�;T
��cfy��k�`	�aB�-�
��U;�"�6'G+��^�d%]���&�".�;��*���#yL�\W�&�I}�[����P������=��ڑ%�T� fg�3��Ξ�Ȯ��JS*����C�.��n�_�	�ۦWl!gu�V�v��G巇��X+�>��U(`\�=tn�)����<�|�ٚ=���ABZ�$s[�Ƞ�w��j�����A
&�=�BX,�)E�yy.2-R�Go9�2��V�����wN�R��b�up�	1�2�L���Ź���g�k�v��v�Z�p(X�MP��I�ΐ�0�i��K6z�Vg���"|@;[��
�����=�1��3�E-��.IH=�A-�(_ii��9��c_z��m���T!�^�CBI�y�a4L���a2�2�z�j�r�iWI� �0�pĪ�ͼ-�Ƨ�߂x��i����6�,���E��g�a�Ԥ���}Ø����|"N�/ssd%�f�`6\E�״����J<��6����#���:ȒN	���
C,�������me��u{��4I"\�)�����h��y����2�c�䋼�O�f�?
�<���D�1�����D��xSt,�v���K*�}��R�~pK�o�*�@�c�@��QQ�ꍄ�[�;�(��|������� �������s�������Ri(�["��.�_�!_��n�uq�T�Ccȝ���9��	G����ƨ�ϒp��jݻ΀�	��p!����M�X�D!�����n�E�1�6�̠=�������}���9�o\���-��ț[����'�?7��̇{�#��i�.�_��K}l2*�u�E?�A%r�'ٿ���2`;?���R��
ĥi���ސ?�.=�A@�\k�����_tk��CQIE����Lg�9 �#��3	��} <�j �̧j��$Ls���0����g��G�ҧ,�Z�[h;����S�p�&�*4~���[X �G��0WL��X�¨�=^��OY{�K���*7�ak�oV�_YIɰp��\='�?�ѣ�.����)5���4��CK֋��x������\qicЇ��̇��������ҋ+,�x������E�j�mB|�[V����)�U^��zsK�F7E)x��$&��^zaЍ�����B�i�d6:-L�(Zm��<5b�r��n�Glzfy~S�K��7wp�S5�gbG���B�o6�E�ޗɏ��uAY<q^fQZ�q���2O��lq+�W�(N��X���А(q�v`7�n��� kB]��a� �^�پx��^���~��4b_��1�	_��$(J03���`�9L"��ӑ�C�[���z{�O�.�f�@�y�D?����;����j�
������G�R
D;�ʩ���"׃5�(�NһZ�Z��w���3yB������+�����G��c���)��i����y�~:U:��A(�I�A0�����s��|m�ҹbUat]��-1��*�^{�Q&s�Š=�ב\)����A�������&m�q�A���Ko�
D>~EL\��P)��)4V1����oOA���$P�6��(_t��U�@����ܩjQ� "�	Qߣ`8�*�*
yݗ�x����v��Ije�^�=B�z��[���)<�D��@F���/�����f��(�i�,�,"��b0� �����h��`0B�#��J�/P�6W�l��}�v"0,r�M��"xj���Ht\e�#͵@���f��-�蝕���܄&�Jt��^s�L`7�z�w8�ť���1U.8�Nq�-��*@���,��� J*��^���<,p�:R4�����*�ٷF�,�D�۫?h�R7Tv�C�E7?��(���|fϐ�x@�tF�èZ�ļ<̹#�$�F��Y=Wb]�_\Q�%�g3ym��ᇗpx�TdU�=`��-��k��F�v��}�8́��G"���ygϾ��^����z�j�$�/)�t�ķw������/�Hc"DfՕ�y聐a[��=��\�t�9�����G��'9`��yb��ƍ�~Q�%�Y+ԾJ�2��h�/���ڄl��.�ƴ�������Z�5�PRr��T�ԩ,����*�+j�{�5X�����HHV���F��`ZS��G��r���A#U �&F�;}QG��Q�K@P�E�g󚯐Ϳ�T�q}�m~26�6�[��3o?7X�E�?��R�_��A�4�}p�1�� *e'���h�EkQ��
��,c�|���Y���$߼��&�;"U��ן�#�R.f�����G��8��/�,��;H	k��և���gJtz�'�!���~��X�]����8�k��"�Tc��r�����w�z+-��䎢2g�m
����ϿN>E���䂽9�1�z��a���c�'i�����3�X��I�.5��M�pc��IWN}�Sd�~b�JD��G��#�,���DX�:����U�=+���B�]��ȷ�o��:lլ\�]��&�\U\�ԩ���[Vu��X/���^��Ϲz9�փ���W@|XDR��W|���踹|J �W/�큪���;;�1��Ƀ�B�$�U��˲R�s�/���B��cL얱 $<�(����:j/U�Ϋ�~.�@tU^P&Y��	'�� 5�-�265<�D�ԟ�����LA�@	_p�$�tV.�7y> �+5����_)�^�P���WN�
{�X]T)\��_-pF�F�ԙ�81`��KR/+����r��N?_���I��9�予z VWJƥ0�^���>�^�g�$|70�)dq�~�ļ@.|�I(���]�U�Ӡ韪�KS�<2�h��a��>�o󃍚hkX"?Di5�;��
G8��M�j�~a�h#/������4ﾉ��~��70A~��(_��꿪�aI���YI����+����e]}�I�_R��!X���I��y����˰�:�0N�	����"�\-�{Oig�;^j�8�����{�%.n${[F����wb�V}���"�_�S�~���В��fƚ-<�t�C���w���w�q� ��6�W۰� �-�o%k��-J���x�����|���i����J��g��`CDN�i�r���z�����	1S�����}�9����]Y̠I^�꿛n(��	V�{V2���7��A����'QnM9�����L�u�	�1m:~@�D?�,b���b	�HC A���t}Qݏ���Q{�����ۑ���&0���oн�x�)���4�勡Ѭ��� m��#�4���Ih�,��0�d�2l��Qo$�-�I\�:X��W��l�,�Mds�TUxҨ�>]B~~�B(�g.	��i��C��I�bKdQ��Dw>8��v4��|2��������]˺G�qB�㸴d[L0��p��7(Rf�5�5����oO~$���Vv�
S��w�\�[1�,�d��W��ڳ��F�qdۍ���q�t.�|�-�D�!�~e��ٙ���iU���M���Q��.��y����������1�]�����]��(������(T��L&#���s�M�����"s�@�z>�g��倫U����ao�@���NF�\},�P��/�"��~�ʧd>Y�Ǹ�����w2��j)��jN�� |��o�� �3ʩԜ��ս~3mJ�Z	-�r�~~�֟քM�%��N/=m��K���	���n@��q���o�J�����dhN�V}AHlF�j����`�adX=9�Zvk�2.�J�����~�9x�apߞ0�:��7m֔����82װ�()�[fM8�V�=Ҹ��"���_��U8�r���������5�LO2GxM5n{,�M�F�XB��� ��xM��=���8���n/�lZ��-��x��=M���R�3,�R��;��ř�`Qd���~�C�6��*��!�\�U��Y��g	��M@�N�,dx@A��k$�n�qn!.J �y��9����1� y�4&Y'<���
��"�dRL�����N��(��8���!E�Bq���gTᱚ,���cj���G@���zΠh�%��p󩮪B��׀?0��R=�4����d�����i3F $�65�~�=+��&�Rc�_��c�G�ː�f���c���c(*������i�U�M Un�!G���m��2��O�Um��U�GZ�$�[=+��y��tǠ��!�>��Fu C�lϨ���Y�����]v�?5p����FA��5hٕ|�ۢu�ԩ
N������i���o��"�E�F�&�~A��h����4k+�qL��ko�?ļT2 �p��!x�5MfϮT���a<elf��L]����5>�;	�Fֹ�툃}_�q@�H}G��Ҡ
s��%�Ɍ�Gة�`��SC�ն�J���NW�(�P�T�s7��Eg�\��.���4�h�ӎ�5F��,�^���;W6�6o��W��Q=^�$��U7Q�����Qp�b��΀uqm����AL!��D�r���fi�I��pk�q���4�hBC� ��Fd�Z�!s�7�S���ٚ�M�p�s����>���;��>V���s�T����P�l��fgB�O�Q����Wߡ~z(,n���8Cy#V[�A�;�6�]Y�Y�Q��z��M���G��������I�9t�O�~�#���l����O�8-s��*��ȉ⧆����$���b�>S-�u��H��
��Y�c lT��E6�A���~�M�=�4��T���Eǎ���;�3EJNK�|A�DEI�t:!�{fU�¯�R������f�֖3:��ntc���W�������$ޫ��k)�8�{�� 1�H�S����j5����%��͠3�9�!��6˧հ�:����,�Mn׭�l]~�ƌG�v$�u!��+ <;t���h���VV|{��+����,5�jm�6�{J�'Lg����3��:8/1�	U���ɝ���;�a`J�k�Sʔ�j)	= ��L�}���q�d(vlD�R�I\�r�?E��p�Gt�8�+�R�IY#�Q;�]���e�\�v
� ����n����1�J��K忳�*X$��SQe{��� #�J�{�B�h y%�j�Ѭut�D����9�?6H�KW^*&<y�d�s ~	��~A��4���n6��}r'<���+���gh"�n�LE�nt�mhƃ��_��%�`�L��~���\�c�,"/<oKtD�FR"C+��Y,��Tum�Z��-��<b��D��u@���Kh�]4=���C�LY���$�g�R���5���Ra�.�۞�P�p�ޮ ��Z`뺿9�jF��#�׺U���>���z�f�M�M@��|=��^�g�KH�}��,�d�M��rW�U#���y6��ڡ�}�����ֵ�AX���b��i�/��qb%4�-��~�����- �n6�kqN؎*��"�V� y�o1y��@}I�嘧���\���eZ|~�gg FV�?�}QZ�ڀh��!N�u�;W�t�X5
K���#����-������M�MQS�أ�>� %4�B�2M瞏��3��[�2���p���
��]c�`���z��j�I����/͵�Cs6M�:89фt����pE����]�V��#(�xF)Y8L~)h���$�LA\�Jv�M�A�̻]�j$!��uʵ-g��l���aۡ������S��o�>�����r�i�P��S!�$�1E�\aht�gm����dKf�յ��]m��㕠2��-V۲1�F��X��Z)� ]V��oqd9;�pc~��p���2�f�
L�W�g�DȻ���٩�B�8N�����x{�z�u����wѮ�y�
�5�#� e���J�C�n�^��&8����y<�I��۶>�q�O����2qm_��f��c���ǀ��/A ��6!���բ�}ۧ�����j��a���1We�:�c�Eҝ���آ��v�J����K��}0xH3�|�ǂX<���PK��T�#�Ű�֑�b!(��_�-���홎M��8u_���� ��ǹ%�#��|����&6��.d����c���8�E��/���غ$���l,c�����cƱv<v�r�-&@M԰�BSN�6}f��[��@!�4fk$F�mIPN�uob����~�8�P�3�Sþ�N��f�V����O��[}�E�P�2�D�4!?Ʋ���6=e�1Dw_7��l<g�xq�P~����D�DB��i;Z,�y���j������Q&BI��dr6����k�%
�6,Ql"ʋN �4ջ�)��O��Y���U���_�U�ݘ`38{�����P��)�ej7Cu���������i��}�Ӝ�]�;zd����E��ݠ�A�K�l|�cQ�M��U��Y���WF����&pkz�yc֧��X����� �h=� ά��Px��J�G<B��^A� �(�����E�@h=���Yy��!؇�L��]C�J�;y�h;�X�mcbh�>+�o��,�<!�.���g��Ӄ^�|���ͰoG�<*����ZI���Qq��V�����}�W��u,��0���?U�2��NT4!�e���d�	?z�+�qhDC���L����Yt9�btG��h�J�c"���sve%;K:�#(�q��@g�U��I��;�՞,�Cmm���E;X��p��!6frs�7��f��+���aK�'%����� ͹�Ѻ��=���K��\��$��tv������A�W�b�L�H"�Ҹ�s~C	�]�T���TS֋���.GZ��P-S�g��+��~eb>q�}�#�,r͆�gԨy\J����a4��#P_+�^(Y�+��m�1���:]��,��E�hN$'\Fx���L���L����X,Y|쟁��!�抵P����TT�6���Qn,DԞ��h�N#����=F��h�K�
��c~�g$p8*#:��RL�	K;1H\IG�y\}F� �4a�g�k����x�@]�m�nϷL�޵$`fe񑾥��0yY�s���K(��ԓ�_�5���ݟ1�bIЦ���T�Jv'�
�z�z�c�t��y	�Z�o�<F��7�Ԓ��"G������b����Ǫ��Q����5�\�t�)�������O�Q�c���}�i��㽈��w}'�1/Z¾Vk�/���8M�O�Y���"�@0Z|��d%?Z����l�Ό��짐�WŇ��AJ�J�୚��qZ/��!�eX��U���@7�ƺwbp���9�����x~�[eF��a�_Hj�;�O�����[[�O5��b#�ϭ2�&�\�f91�g�;H�;A�t�ѨS-u[�&�Z_�\D������"�R�c���y�>�*�NR����"��]&I��we���	A+w�n�/_*�'%���k��ɘ��c��Uu�_�.�ȋC�����Hu�c:��;hR�耘Ve�&|�/v�.�C�[��Χؾ��|K0����b�J�	^l�h��h��g��.._l��S�-�k���R�f!����ʹm�&{�Ј_�վ�˳���-��,C���\�V"ibdA>`�>�t�B��a������+�Ăv<���陸��cI�����@���QNp�dq�]�������zѾ���Ժ�*�����_��>��M7��X\�/������{R���;D�<[���+�H&O_$/I�pI�c����@\H{��|���z5��8/��{�#���X������X�3'$UR������������1�鋆6
�,2�c��T4kN�"����$GC,x�k�����)��f|"p����5�[s���	.�?d ��U~a�>@A�=O�D L���xT網��>JH�]9�+�V�}SHw�����Qa H�k����
��3�Ukur�@���a~K"u8��"�.�䱔О��Ynb�EѐԲ�B�c��;MJow�Z�{0��p(��kO7�H�<ݥ� n�r-:#����$��HU2�y��H�� ��a�%s�\���em��3�uM�1���{��A�D��$��(��^����w�
)�X~����]��!_3h=�B��w��J��X.R��0u5��񿌰&t�-�����_�+��~�ܝ���J��U��������-+��[�l��k-�L�:X��z}��7���Z�э���G��u��-�1!���<�y`ў��J���h6˓��l��U�=p�N����7?����\���yZ�j�}?k���9z�P�FB���� =��_�9�U��`����u �˿��m����탌}���+�BZ'�F���-�1p�w3i_5��у�&�mL�|C�普B|PK#[��n%���XQ�+2��\4:K7��V����?]��pJ�x�bZu�!k�7 q�3�J����^v�]#n�"ڰ4�dC�:�d-}M�[We�y�����j�5̌��b��ɞ�-^%}(���E��f�۴��K���j+�6�fY����=@	^'	}�V�eg��ucTN�/z6�W�p�w��$�}{�el�֨]��_L�����<�-'����v��B%��'Bb��S+����~���^�E->@Q��b��O�Ⱦr� �Q������X��b���K^��i#a4SW��
�d��I)��4�j�_f�691W����\W��h1��#�7��5�z(�pz��<�>:�Q�2��m!$XpI�cRa����\�֌p�\��ǌ޸��/v�d#ߎ�dک�x���1u�:�G���?VƵ��q�	�\	�WRy� KE��)����O�kOf$���C�i�Ȗz���9ݡ��ȃ�%#\i`�K�*x6p$G˚ل�U����[z4����z�}��(B]�NQ���ݓ���G�+r��=G;?�K�E}�5���"0s>��Pi\����Ɉq7��C�Ӿ�E���D����1$�}
�bEeO�=@q��=Zy�#��$A�Jήk��]i�B3�q	ˍ�k��o�,O�5���< �_�S�M�H��=c�RD�gZ
����Sa�@�u~�w�����]�:���=�r�9��Y�.�{���O��d6B�%�^k6�B���B9jQ�9��Q_1�"{Q2n]m����*t(�ɭg(E �ȉ�|�/Y��M��'���%���k��\2�2�D��~T�o`�ӻ�����2��9�I0d�K����U�R�+*��W�j�k*)�\M�ԛ'ڋ�6ڔ��BB̬�6���m��ަԐ9�5�=�
�3�v�F��u��,ݪ	����[4I�8����(D;��f��{���^��z�ſ*�sD8l���L>"4�0�͖�w-���o��Ǖ�\�s%���UA&�<�4�	�LÑ0^ޖ>���`���}�;/]L��e5��W�չ�S���_��s��H[��E+���[�ݩo�2Mb\u�	����=La8����V�tG���96�?<P�qtI�A0��i@����*75A�g����j0Z(G�tH�Dr�o�y�˘�Z���_g�\GV�����J���|��j�> �EH�v[� D9E�����CQN�JZ�3��Ĳ��D��n	���ϯ�X��#zD����[K"f�;�Eɦv>^���֑��K)P����V�$q>U���ڑ�����A}�e�H�n3��U��.'���El�]:�_���/׫���)ή5-�֙��
�*>�WҨ�6��Jt<��u��	�\�1z|g��ވ��GW+����!����CPF��l[�ʨ�,��ba�כ�q^i��jy{U"��-�JU�H���$�_�j1�<p��w��e�n'��0��1vb~�	E�+�;�n޵�F\��ard$\�p��;~B��k�g ��x����^���Pм"� ������o� >d��m�$9����>���m�������)��:��-Dw�W- CtJN�ڨF���\���Ӟ���y�]q������0��5_	�9�<�~@��:�����3�+*KHD�a���^�̝��d�fxur๝��6[�W��kn�9�K?��0�]/_4v@���{%:��*3���i��ʦќ�cΈ�O���LI
Q��zu)[X��	U�eg�%*Eo�?�k�y��&�B����J�މ��ŏ��9�Zb��X�z�"*��(�{����X7X�O��灥k��#���"�#nmJ� ��N�vD�`�Uߧ����О+������(�l�wXvC�-!��GT2�[RS<��r��Flmd���<�1�C���&?#Z��?w� ev�_z+RBJ���~}���vƵMåX��_1!^z�P�}�� ��%�V^��j��2#�o�	qL�%i���*V�f=y?>�T�+�7;�}K����.�@w�q��t��wA�>&K����0���pd�%}]�e
=Rk#���~��?�|c%9՜3�>X��2�ݢ���)��긺�l9Na��ʃHk���`V-��e&�(\��oF�Tb珖�򷍵{�j�L��kqC�9�*q�~ w������{�s�F̻Jq�L�#%���b)����s��%��-/�pS�ތ7YK�3�o{��&xZ+��ߏ���$�yA8{Ć۰�����g�l��7�o��gM7}`%��T2��e�E�6�qX���:��Ky��.²s��#�-�� y�C�La���w���nURlb�:+��n:ʔc59A	5����K��$='��1jI퇭�"t�`# �df� t����QEz��d��A{�I@8���@����Y\��
&읣��s�%L����X#s������bG���Bfzv�;-a4i�K�B�ҟD��7Jm=�b]7�H��7��Z�������S��;�w�8�X��!�#2K� t:������t�U=o� ��m�'o5"�ܹ�y��I(�S�("�D:Z��y��%E㼷�ئ�[�*DE�m5�/θ�I�+o�=e!��j=�|�ӌr��2���ҕN��2���Ǉ��d>�5���Y'3K�Zb���e��A�'��}H��ia	xH*SH�g�|�:Me����Z����EfI��4l��97qǏ�z)=ic��m��90y���#{�H2�>M3cEO��&�v����̛�%�\,Z��֮Z�Q��w�UkW��n��#�g��"j��kL���!lҧ�z�A���5��:ɩ�"Om
���(�(�S؀K�ZU�K���䡭�ⅿ���-j�X�Tg�֯m0�ne;��"F��w� /ǣ��A@�x�1���P���{ɘP��T��G"h��d������X�i}���lo���fMe���;��$dxE>�pϹf�<�"��d�Y�GN	"$w���Y��II*0��D'~Г��ާÔj-UA<�8y�����Ty�@)��v�����x����7sSo�&��nz����}�&�;X'�ۼ��i��%��yazp���u_DŉzX��`�x��/^,��o�i�폵�Nb6���s���M-x5��,��۪�PÉ_F�2a��;j��J�釚����~Ռ(7z��ݏ򋇌L+�F@�ߟl|���%�5�|�[�p�U�=2H0�U3P^��Y�8�<�ft`�$�;|R_��w}�?X�~��^9|(w�C���X�1��:O��1�����n��r�Ex :.�ċ�8��m��f��u�����9K�Ǫ�_���i��W�%�( ���]`:�_�_n�4|b��q�mR�;�V��6:�%�/�A}�]g;��N� 2��3&kuT7��m��/t�^Wk�T�tCn�!M�n/'	��K��i�H�d7�+�t�ׅ-��N:U���Li��j���[�oT�C�1��p��U���)�8j>3�}������!�)���iO�ȇs��,P
DUH�O,�gq��(�`�c�-^_k'������v��H�W2�đ
���v���p��)|
�5u�x��k�i�������⑻�%t�z��շ,��F�������B�5�`�?E͊����
�3�[���sHS$�CH1����j���p�m^+��oH^νs�*�ds;(���|?k	�g�������wi���@V�,��4��z��I��������c�Bښt b�a�ϣ�.F�s���\3jIf��m��&�p\Df��(����#���9���$.���g����Y�̡��r��AN�t�0fh��r2��P��}�F��Ð�ˀVC�=�^%�qB6
y.��������/��C��1��t��-c���Q��(B��$LYiH��}��`�=ڹ���irTv́�����YZ��atȆy'x�uY���K|e���hA����s�TI
��Ch���$ċ�ǒ�V�9A-�}� .b�Є�FA��M�\��؜�4Ҷ�'�Q�x���ʧ���r ���_��wT�Yw%�m���Uڻ ��G>�`��XH�Q�L������������nri��I� �-��8e�nR�����
%��%�s#��h��JW��X��'�}n�Nk��E�q���5/��0"?��0�u��"�iI�S�����iۄ��׆|���tF[~t�!l��!nK׋�MhC8�r�ֱ]ݻ����9����r/HǛJL(�'�D�l:�O<m �X���F�0���{�3� =�Q̔/����a���z:y����l���Ez:���(x`)�)P���UY�(�i��,Q�f��QP%����zcc����4_+"���H�5��
����9��UP~�-�7r眍	����_0�A>d=ד��-do@�2!X�D8ސ�d4����I��͜�7��;s��|P��qB��g�D���F0��sLٔv����kt ԴrS�󒄮m������Ǯ.�)TՊ(��kE�����7f�����|�-b�o�!����"�������E�C��M�c #?���4��nt�z��x��4����q�f4#"��~V1��G���I�oq�6!�	l����|g�k:Rb!�%�D��� ]0�Nn�AYa���Q�f/|0�T��qN�i�hd �n�3̗�2�"��[���h28���J!����O�x���u�n�9�Fc�o��J��c|ڍ������&Ź$O�a��t!�	��8k���}i9��v�Ë�{�wV�4��-(���=��J^�
��ֿg�kY&Q=�J�h�̓t��/�2��d�љ\d~�L^.��GS㜧��]j�X����Y#���v���&�O�������A1�AݠZ.�����W�5,/[� ��GM�2a����;q;6�M5�X.6�q�#�``T�O�X�U����Ԁ3D�834��X����~E�d�P��O�lv��fp��mg�p��j�%�b=�~�� x������'�M�-�<�7��mc��2�)^s�l1|n���:�	�%�`��]�t�W��w�x.���RN:Oӄ�o�F�+mf� �G6�3?����<%cƄ����P���8�"H�z����?��Gh���0ϙW�@��o�vl����i��� �O/���3�C%�����'L��@�F"��)��}$Ŏ�p��J��<�c�wI���W�g3���~x�{v��8<�G���f]�2��j�\E{1,M��G|љb�j��R>�d17�fv�4�QP@�+��'�xJ��<�C�˩��eY��/B,1�mqX^!�k���oY�q�T�)=y3D��w��0} EA�q�4�2����$��$	Ch�����1G>���a��>)R�4�{Z�����#�h/���i�K��n�>�G�� ����|59�r�3	Q,lOPY�^d�Pڠ�?���W�x��N�3Ix���=�
MU��v�E4<� �{��lĺs�C?�<�۠ۚX�+��x������|�6�,3�X����E~�HW =�N�/u�'��ٮP6�9��l��*
�"2���hq���ơ��qzDː�����#��|`�ēd�5��g�� ��	�5��A: �`fd 0�oG!Q���Дj�$d�U�룿b1U ��BEy�)4�/J?{ET��b,�ޥ�Y��M�U[���r�;k 	#ȉ�#��UB��Ѝh���`��EF�}Z�4�]�<� +�Zќ:G�lQ'��=I���Ő��1q%���9��	�݄�/9$�Cb�K���柆ؔG'ݢ\��q!�Wi q���{Gm��- ���� �o����l2f`��e�l�#Ui��W�*tY݊��p+��w:�����_�٭p�����L{9`A��t�fC�"˧5��5U�ηY �����Yd�&��:� .Z����ꑔU��I� N5��M^�z05,fU��Y�"�ro�RHw�La�,�-;��Œ�`$�i�u����uu�]�ΟϨ4v�ca\_��>4Dvm�D@.��H'p�=ɇ��;%��j��7g~Ƣ�g3���bd�_�
�S�Ku2���F@C�F�1���]�D�������x��8���>?��"LD��Q4}�d%�l�������YJj��Hv]�bh�H��܇e��z��ְBe���P:&�'�fC��.$piUMm3=:~�����A����>��Ias��3�%-9�ݽx�"����d�G�����3���vD�n��>"�����x��b�$Q�Zch	/(����Ba��p�X"�\���E�j���w#N����e��^�C������.{��=�D� z��!	��R��J�"߄b�d�Տ(���2~W����M��u��$g�=����^�\�-G�X"hnD��Af�6*O�<��dH�%�<m�+ԂG�ĕ���x ���>���ݣI$#$�-�m{,�܍V@����"��y����t��Aa�x֢��*>�������~�n%d	�&���T��qI��Ҷp����}K�|R�(ؒH2�l���D���J��0��ҫ��P��T���J�@g,�3�d}�b?!<���&�L��%���}2|%Ok�ab�Յ>�b8�lͤ��'�U} ӳw�����Iԟg��������+��Ak��l-u���f�¼>>�F� G[
UZ� ת��j[�U!-�e�ɺ���"@$��Cy@�޼�xU��(ٸ�x��g椗t��Η"�����K��x/�BL�ӹr@ ��lE |��7����?�?F��P%Y� 7���A]Yɼ����_���|�����F��y"��)ا͋�8�	7��B��	�^�qf�^/�F��U�It0:�ߡn�)��p���f"z�9�8s��86jG\q*�����YSJ��#�"�Q������U�40��`��R��d�����	�,��T���_�V ��wy�g5�y��x~tI�S�� ���M��6F����2�GlEg�%�{5�t/N�1gP~3���B~���5#iά.l'�2�J(C�8o�3�C���9���+0X�{��C��yw��P����[d ����׀4���{Y!�I@p�p�%��qȏ�=+&�Ti��^C�d~� Up�}|2?�g3�+���~Eن�V�ԥ�J̚��� M���:��?�+�'�{�?�JC�\�P�j��O���ؠsx�H�%a#�n��D�ʢ��	�e�H��BN���N���M��$ѩ�����w�t������A��>8��#+�v�)c�5�LĒXc������ �W!/�"z���hy�&�=Q�lj\���0f����r��k����,���+���?���ǖ�.ӽ��@�#��!�<�(���5'��'Ce��˻�K�1�ϡ}M�+����b��M���wu��Q�����Z��.+C��9����\i���[В��V����7&��j	(�0���n���/b#V9�~��	�b�n��]�+��Y��Dϖ�EA�q}�=���Wba��ѣur�
h�#5�9�͝��Y�>�7��xn*n��<�_���qjW���9�7����N7�ˉ�o;4)� ��i�[́�Z�^�!�
#���1��o!2s<�#2�"B��q)p�js��wG���M9J�/:��[i���^���d���`��.��0�UÉ(�2�v�����;
������q{�`gLЀ�6b�Y=@��!8��"�|����]��K*��6�v��
�6&;qQ�cL)єꀭ,_���Ad`7lK������L�S�3����������.��ˤ1 5ɢw|���D��_�\5���8w���u
��!zu�ɁD�M���->�b�#c&�ZX�:�<��� ;W��6�Ž�'��q����| �B�R,�0V�8�OK��ya��~U)�L���C��M`){�*� �33�h�[���]L�Vz�=�g����mQ��6(SA����p"�J��ǳ1��\��[�9R����*@e�*���Ǐ΢@�L����
�2����i��8�� r��T@gp���'��"��$��
����� �;IO��	P����W����+	�vi�D�3��|h�X#�����5UL,�k�_0yG[���b~�i�}���s�Š����Hp�`:En�Q�& �Qu���y��RO:
o���-Np?�OT�1R+���<���O)I�t	g������̕JDR��z����d���~w-/5�����G���$
��V�8ױ�^��U_����l@PIf�'��+����a�!S��ֆC�gh���A�U�N�������Ꮆ���D�����ՙ"��8��n�c��{+.�D�f˜ŏ��3����p(;�M+�2L2��p��;-6�2S`K���ZR�f2�N�ЧG�z1[�js7C�ͯ�^�8U0.u��� [�_�X�1��REШ$�{S[��'�RM�j����|7#�����צ�CD/'P�$�t�}���)���K��{���0iB�LWxΣ��@���D���*�L3rYl�E�Sa����p��X������E��<r�����^���Z�D��E����^���yڞ��nI���ϼk�5��&�С�+�G���0JVU-����ұ��
�� �%�.^ D\�J��������Zdb��ml`�iG�E�#";E����!�r��5.P���ҫ?�m~�[��]zۺ�!����F�k����vc�v+�Ri���;PY�̽��'����䬿�:�!2m���}�����:(�D����fFB�a����R�4E/�@���ly��0B}V�Rm\�g���k!w�#�A�=R[C�(�{-�yj�V�gQ7�M-)��f9�P�`S\�^�t�UOp���LP�G/��*�x3j�Ҕ��v={�s;`�Z��2Fy�/�� ���W��Uǫ=��/�9^�?}�@��{��2�qEt�o�L�a���W��CR9�������{:��s�<s wq���<�4������-�7�\�C΅��8�w�"��X�#�.��{�u
�@'�j>t�<���F�~y'��{��	KƗ6a�+��
g�f6�7�2�V	y���*��I�8
f��3~�S+��;ABZ�}�*���'<�_��\Tr&�cy�<���xi���f���� h�{�n��b�w�b���ש�s@5dZ��@(G�,��j���2�� �R�ۡ��WҴ���N���-)�9{&R:���1u� ��A�-՘p���L���g%�6`�.[9���k����!}���b���(�&t�t3��q��n(�Y�����w#'t�	���lR���N{g��7�P�lg3>���A��_�]lj��t?���2�L�x�]�G��l����$�:)	���,�28�H]�A��Ί�oIQl$o�.,�ݼ�,<�
�����XP����������}�`99�p��ǻ^��92��xP|	,�4wI�RɆ��+�KZ0��]Ѯ�I��d_�"3����W��]{�m�t���"��B�q���?J��zv��!�C�=N]A�3?1���v�7h�3ik��X�)zz	��{��c �D����W��:�{�d���N5B�0!�^�ѓ�4�m2N��y���h{�h�4�� Y�Q��>K���v������
F$&����$����u��(�=��;��.�􊝬�,8%E��"���Ά}@\t�y
	.�z���a�%ԑ7۪�
��Jgn��L.�ٟ��X�TAy��	��ܮ8F�O��NW|�и����1�����8y�g�Ǹ��r�tY��}b��=Ꮦe���$rS��F)
+��V��<K��%K��d� !z�60�ߢ|R^?yo�y�#w9����
p�)�?�0���=i>nb�  �g�Pl��l\�v��X�`[e�9Ct#=�K��\R$�����|�Q0�	�S�$n�q�NL��8��L����S D��"�&����E�u�9���7��XT��Ag$�h�}T��˷�ez��>e�W�!e8�|?��I��yM<Vkm����2t��g���`ak_�ށ>�[6B�O�
˾�i�!�+{�#[W4��Ss0�H˳�� AUG�:����Wl�#�/��Bw��u�K��ˌ�n��r��DMU�N�#��7Yׁ�������{_hM�d����p��.��W2��s'�a7)	x׳V�{�$3C](���>�t@>4�r�F��1�`ۏ�?J�O�dv���.z� Qw���n8���m�J+�P�=����1z�bi�� ���S� _�d��vQ*�ڪp=��7��uط�o\(.ɳ�]֘{�2S"���А��+aO���3E���:��2����(p��PgdG�%��j3���m�G���:���x,�F�[g6�]�:`���8s��ɬ��B0������+��A�4��x�(��|U�f<F���7�+�� ���s�^��@a�f��`J$����f �
aXW��.�,�%yxP���(F���U���3�����!O[�*Hf�͒��/��m�!�3[��]�Y������H/�	ec�&_�r��A��O߲�٢k^�@���fԎ�5��<����(n{��ȧ�ra��]$��q����\R�(�����L�����l��<YX�_h~�G��x��H=Le�f���s�1<�w�Zq���!n�l8��v���f1O���X�jݕ�8݌��]Qp���T��7�bkp]]Ȩ׺�@�s��-i9Y�_Ue�es�2�l)r/kC�\���IX�1y	_Vm��\��S��V�j~v�f�x4����-0&�Q��vy�{Xj��"s������j��$���������E`��-G͏)����Rˮ:�n<�]����ڰؑgn)iLe�\z�C̲��H�ř/ 6�:1�G�Smz~�-��:SKn�f�j���,S�����Y�>�0�Pn������QZA	%] .ؼ�e�����vVK`-
 ��*)��2�DZ�r��9@I�ɜY{�k�NT�t݉Y�i^�j���0�04�4���v���	���7�^ ����o��4�i��|���/��ڲ�&<����[����J�|�8trǂ&�&����wh��Lz�J'NF���>A׽��	��k~��|B��lEJۏFp/���I[\��6��E)���K݁A;F�!��\ǔ��@~��6w&��c�z ��-�tŮ�ؽk�6$@J��̈��%��sn��{e�'�2��Tr9��D���6����X7at�v�W�����
�K~�Of���ܥ�������i�1�[�g`J�e����T���^���aV��j��/?C9��Sb������ܨۂK)�0{�ϝ[�{�K@������5(��b�u��}"��X�[|+૳ӄF��
�Y��,�'.���Q����$����������2�c�.�]��u:���m��'��Vw~V�M(�M�:}:G��&7@P���}|�D��Dظ��������A�4���Iu�c2岷�Px�J�
��o	�=4��bS(��S�[�%���*#aN�=\�k0��}]7B����T�d�1?p���P�� �3��в����Y��A��OV!���I*���O��V��z1������B� ��`��^�̠�p�.��E����'���3���hD���E�{k`}�i��z|Q��sԭ�/��"���蘻�@��C����u��̅7��%]e�=��l]�;��IyZ�'�o�Q�����1�3E$D��=?��* JJM9�v�آ�bS��i�� t���tJ,�z�㨎$�z�ciW�@��Re�%���oRI����c��ɷV�wڇi?j���,����cnax8��^L�-������k�q��=;)��o��b�1O������G�\SQ���_U��7˱QT���G�: �ը�H���c�̆��aT���cZ��Ҹ����ӎ�-�b�)��:�Nb{�.����<ci���E�FK��|׬\���a��˯s}����΁]&t��/������s��v�c;E|UQ�P���dJ�ҡs�L`�B�la�E�ӣeĈF�v��jPD.#���0��p���!lF�R� ���j�U�m*Q_���
&pc�A�z��rEb
��6$E����V��
M�>�
�/�<gۄ�}~��t^�9��<b̑�:[6ۨ:(���c�X�c��)�Q�.��0��deٞ�guw��v�Z�N�D�3���,0�|���k&D��O�|!�%_�`�5�-@���%<�|�|2]�r�=|���W�pQ&���?&Rş��Ӭ6z�W�վ±).�l�ФZ��}G���Ğ`���KlR�Ӽ�H�"����?U���?����:=g�K�TD{�;����ENKv�N�#�Q[[9w���}�E(����h��Sk����j�%��hS�A����6i�U����/s2���(�������J�i���t�;�j��K���f T4��jrr��
#��MP�c�f��~��A
f)���2^��|�˟W�T�v��ε��)��"���u�
^K�~��������M��bh����(�4l���"��(��P���^�ӵ��2��%,��4����A�y��y�󪮪f�lZc1T7�xc�� s7!>��0N	=���5�2u�F���u��t*���K��o��,��
m2*�Tc�>�AWz&[v��j�!����`��*��Ĥ�Bs4>�"����cAb�Fmlx4�>ě�
̶�ϧ`�!Ţ�i��$f�f2�]�G�8"�|�ʆ�дb?��9�䤨7�\�� $����x���jԐ,���5����	��:�C��Cg�I����YuPK,[��y����Ee�{�l�P#� &���w�Vf�A��?Y��$�T�eB��6e��>qe��")�鈴�tu^��1��ó�Q�DN�����0
����+�r����²n� 5���B��%@(�xe�#�ЇJ�e��� (fn��J���a�Py��sZJ!D�u�A�d:�Q"�[S�}&����pa�\Io۞$kO��do���FW{�K��^�!�\c�o��ٞ$#���+��ݧ�J�KS��'F6�m?a�8������� ����U�	�
w��� ������ 3#H�c9�j+�je��H�A�G]�x����^p����.ӄb�7/;�{����ԕPƘt�f�S�3�	9>h�Ӱ�i�>S/D�a���ʩKʛnφ:Du���;�>%��g�k�� ���v)�mQT_���]#�k��e9�ցp�
~Fk��e��0������ۺ�4V�:�F���X��z��T�Z!�') �5#'F�7D�t�] v�O�`"�O?�[�14�86�3��]�Z [��l�i�A�-%v�bwf6ѯ���%�D���	�w���&<j�9����ƴQ�O�zH���W���yB�PN�r.a��~v�x�(�g�٩?�Z��g�"�U���,L���x ��:���З�\����N�����2���^����e���&VÈ��㵷;͆��s`$g�]_$&J�p�i�L|���u/?ұ�̎G�P�%��P��:���d4ڜ[�ĞW��ƁN ��	Z�[�[]
X��i��Lʟ�,�N��J�莛��GQ�o��οe/�
b��I��S^/��)���R�Z{��u��#EI =D����;�5V
~�k��I�\.�I�/w�m�dvc#MbMnzyE��Bqx4�����!pӎ�2Q["��E�k���B��$��#g��OF��:Z�����%��e�%:�:�[Wa�����F����7hGH;I�F��zD���p�c�fƄ|�t#��b���u-<gQ�Y��6j4��l�r��Y~�Z�>��^�}�%�1�e������F���a������}j�����bq'M�a��-���F�q��	�I�xy����q�(���4-� �;D��Ae�Q�U_e�\����З2��9ս��<׌p�n�t,#������m(UDb���r�&B֓?��Y���D(rc����#�ݻ�������:��u���7ea1�2��h�W�����Zf���$���l΅�T����]�/�U7@y���L�Q!�ĂJ����P�j�471�?<;��9�GkS�p�He���5;y�Y�{_�DV ��
�)��z�T�m��t39�_�J�vy�����$'j��98�Qb���l��H�w�߳&u�{���]ojq�*��+�N���EU���佬v�"[�Aa�'����/H�K9O�}�Ct�6�Q���7��[H�$�A�@1�W�^�5k0�x�.Tz?Iɸ�m�L����CeK�	����_���A�?��Z���fD�^0Θ��!��R�zG!͹j?��2��8�AE�U�C��!T�����1YF��ہ���Z&w~��f��H(]�^��<�q!*����e�:Qw��v
qS�=��������l7�kB�Y&wvJ�M���`��,��k�h�>�
��{�G�vE8��~2ࣜn�����B�Vc�jz�S�aQwf�V�ǉ����G�6��\����K熫��7^�O^If��<��S��8K��|�H�8�5�1�Q`Q��,��n:���$7�㨁���� J��*����γ�mߋ���0����Uo�K�� ���j2�Ɵ�w�#f��!�#�mK������PХ�|x�Z���}�����"a��;��Oa3��X��o6�Jko�;��,@���d��FV�8F���f�o��(��I���Mz"`�A�!�[&,��ދ��К�O���Q����VnfƇX|�����������HS�@S^>7��f����J�C�ϖ
�$I���c�͇G/A�Qu�h����ٟ�p����],I22�M����]"M
�)}h����FVU���s� j��{����:6���eb��G���Z��0�f�R^�!�>�^�1�lpVP�ηp�{m����SR4�x�4��6<��<]�L%L:V�;�2b��K��5.���)��YY@r��}����D����C����0D�| �,<�$�K�+kvw6�U�UdV,��R�Փ\E�6�Nޗ�3�9�oƬ	ruw�F^1���Cy�F~��gY���H��7� �� �|4��x�����,�*�VI��P��X�i$l(<�����⸃������uC��9�&�$T��l���/���N����� R�!�Ǘ@��4#^���'sc^<���A�A3�	��@� �d��)��*����:Q�2��{�+�n���4�����h�TgO$��}�n�hv� �>iq��{R,SK�?�*,�sDÈY�๜���V�ѵ�O�l�v�g��p���-Pm��M
�7�����]�4�V����9���������g6]�����`W�
��-���tG|oU�p.	�}t�KV�W��B�ʑ�ߣ-�z�=F�6�k� yz�R�H&��0#�����r��[չ�Ⱥ -l��f�N�ǰKm%�A��4��Z@Z�J����t��M�]tc�6Kd��݂�w����0���;@
�_n�%`qm���C6��2'
����%�P�O�]�=}V��/���m���(��p  ���ߵa縷ן|ܕ��E�Y1�iXs+2&Q�$~�khy�<m��͙:��c����T�B� ��%r�Z&d(���*���3wI:*�Is%�f�� ��}H)0�{��{��nՀrQ�vwvc��i,<"�w��!p#5>��~�z�2�w @�|+����"-��_P.��B�(��P�#�O�_a���G�nl��:_��r�媓�*I"�+;v���ߓ�9�,��L��i�S�m��M�^��v��C)���ɭ�&�e]�͂k+ɛ?�9��$~�)����i�c->��b��d��7�#k�,Y(2��J��9y�[4Ԫc� [34��<�M2�p�����ſ��������~����y�k�m���#b�r�������30]T��s���D���Q��K4�l%�ا�I��v��)v8+��Q��\�]�z���ܩLA�����
Ў|{y����EN�?��QьB�Q�$�b����'�a�NP�d�æ�mZqf��-� ĥ�o[1]��/����uYٗ���MӘ��FgV��I� R�	9�Aۧi�$	�/�f����L�k�^�;y欉�^u�|�`k�pEԂs�]�������3�)C�v�H�Kp#��&�Қ9�2N�İ-�2�h�;�ݵ&0���k�1'OB���y{�@ו���\1M��:/ؘ�"����}�T��}/��[��]�6�V�_�u2����m�D��f�R�����-�(�m���?%�(qb���gZ��$6�H7�4��=�f0��~�k(w��3T�ԝ�=	u� ����0;i����/F�4M���J�H �,���P��]����s������ 9���t��87�1&�l0�*).D�x4�V�ل��X�GAf�aeeuEK8�������Hj����2��;�$�'|�J2C�K����<Z���@3MɁo悽�Y���T,o����OU���:���l�ב��aL8���zxjmu�s&�B�e%wi,��}��������ݴ��%l卛�3 ]��vŐ�b*$�.۹���Ѫ��^*�����!H]���1�����kxL+jf�]S}�Y���!��=h���V��`�F�K�R{���\Z�xAZ��޺mHb��%xo1��8qI���g-�����JFx�x�T b���x��|y��S�?Ņ���A������#a�ԐC��Kv)�+���-��ݥ���{v�`��8��hQ����4�7Uȏ�:��lKok?�æ�k~�a��[O%���������D�i��Z��[[����}��.��=;��4�5����3�-km{_�Vy�{Ph۹�|�>�gGq�,�6��@Zg��p�ۖ社X����_�P`&�d>�eK2�m����w��v��v��N�.E�WWV7R���Ց@�ؼ�x��L�Ҵ ް��)�z���\��,we����u��}q�l���eO��������.S���A����^壹�����`�U	9��q�Z,י7Ym�mn�V�����k�����ׂsNt7{Ш%$���.�����m&�+�S_f��Vx���{l�R2H��? �� '���G�3�N=�?Gh�5�qo�2p^V]e�2�"�Ybգ堭&����]D�@���&08�U�鼇�xg}���;�`̔ ��7�a���U���Q
��|��a0t���tGj1�u�����%�$!m�K��Tww�1��� m	Bꐊ���j��;�xX��h��1��+�-�1N,آW��[+PW��J�&j� <B�I�%�����>C:/�'��BƬ	�%����������?��R���'b�8XH�rʄ-��㛳5F�Ru��ٽ��tf$����'#�F�c�$�G��a�m���8$|ĳN�O�6lJ!W��V�9����ua�`�� �4�诃�Zj�	��6@huz����b�k�]weG����"�x�N��MQF�r>���e�WN��,�@���`�	Nv��gC��(��K���m��� �k&�����񣡻���g��/�.0�w�	�N�� ��`|�`����k�S鬼K��W�G5[���R���|)��a��KR"vο=U�rޮ	���N���!£�	xL����Kʨ�ȗW#���a$d"Y�����0(��J��U--;{�엮�h�>ə���yp��4�����O��������nX,i@TU�wm`��I<m�< �h�l���x��kôS�ބ\��K/[g��p',Xb� S�jQ4�{�/�C�'�VM���O�i��R8Ǵ�ss�{mΈo�(�x�������(��çk[z�8�`���u9�Zf�lF�l�ڕ��
� Y�������C�EB��\�-QkW�ZK7��7L��ё����\1��n�u;��/��Y�΄��A���C�qCA�����+��po�,E���ͺ�MǏ �۴�5�%'��ޯ�3V�	�\ר�?L3�Ni�F�f��\ԒTI�}X��k�2�ʬ��ae�N>ȮT]\-�z�:5�>1�ٯC�Ip
�P	�GS��׽ Ԗ�ЭA ���WQdS���`�
�}��z��G���c��^�!��;���0�֓^�$�X.
(����~���Z����}� �(�w>�̈8\T��}~!4�\��<[�E�ˣn%u�ŰFo��5��	���eR�_L�ޝ=,q�J�A������-�*�p�b�{k?�W\m~{بha��b� ?��@��u�g�d���&T��x�=i�c��>WԽG��� �	�:b9>UX !�O��8�8�_%�6�{�|!,d����� t��H]+�t��n�����˚�)��Vr�������Mc��m�d<!ޖ�������M���Z������[^�7���i#//�S��T���a=����n���1��G`����ӝ���ԯt4f����b���R�)���:c[_�T*�t�����ͩ���ceJ$��j6�R��_ B��G�8��j���&��[s�Yd3Q_&?��M�"���\^2E�]�������`T_��rN��E^\|�W�Gw�/aq�&q�nF�ƾ��g��'�v�p�p5�M]�߶��f9IC���(=����4K��L�1� �)m��띪���@�,|؎�v�&�v;�?�(�ܸd��yF�DTC�4V��}����ei�,,���pC-	l!ėY���T��ަ�~��m�a�Gn���_�e��6awS��k����r��,�����n���_�����q��C{��-2���8��
��9D=#�1���#��Ms�/>�.�c��E(�NHZ�1��,p�z�aQ��{v7R�,��8�Ӂ�b�C$�u�l��a����j�T�&��K��b̃�Y�1gk;�W_�#�2���+Ny&�eG��]E,, V���?�)���ìZ�*90��Z �;U���hU��"���3r�L}��T�J$#<������h� iY��^82ꇁX�����!�+?�������ƅ^�u	sg�����)\�ج��R��3���d?�J-MH6L4���}��E\E����_��S؍}�����7tZȅ���N �}��2.X��G�Q�E��o��R,�*�K�#����-Y/�2�Eۮ	���;�C��)˱p$�/Z�����P�q-6AA�dť��ؔ��jv�[e����φc2�߼����E/�+��զ�+0g:[y|ʧ,�,0�҆{�T�S���!��E�U�
0�4��[8�(����2� C����\��.��Pꉿ�9TO!���"�΍;Wx>IΪ�]r�,=��W�WA���_���[~����<����#�6d��&����B��KuX�S-�_O&�N2L�k��/�h�g���Ki?w�0m����Ij���1y���O��:v�#�|��ȬtV�Rk3��S�\��ۨ)�e�,w~zd�˗X`8����ј���# b�i4����bJ)ڧ�~�Ѽ���g�J��3����j���f ��̳�y!^�՝�`����,�̻��Ԑm=*I���e
�Ϧ�2���.�s�gs��d�6��`�v\FW��T�`p)"⫇�*Oï%�tW����0���)w��z���9�����Eǹ^��p���7ĸ���Κ6�{5�O]N����O�U�<bht9"_�*鱹%c:��x*�a�jD���l��~V�����}!i 1��	�L��PZ��2����]�/)����T��p�\.T�2翓��L.د��UW�2c>U��<4q?g������壭���C|�
>�S�=�Zp�Rx8X�}*EI�hl�5�������,��Y�I���l�*gF�L�/�'~����i�L�.�׾�b�\�[�H�+4)�%b��w����d>>Т���"Y�љ��@�#�SZ�2��@π( ҉瘽�>��)!u��[��	r.�gB��x��YG�Z�s�AM�K�z�����ua�l��c��3��O��u�fK�q����Z-��<Q{a�����)�>�-���bp{[�=�8<�a�+�3��}lZB7ּ��dm������R&������'B[����� ��C���'>�������e%�l�QV|�?��<-W�@�h�?7*�%��\e��
������d(�l��MVP�*�S	w�#S��.(�Ƃ�6Z�/ө��/�G+y_5ս���3�
��O�?1�L����$�h�^�@�kѺ�L�������H�%�V���`�7Q)��@�o��/�K��UּJ�BT�͖�ھ��Qǌ�ֵ#|�/Y���0_6^4M�
2��w�f�|U$��tw�	�����Ǉ�D�z+���G��P�vV�R�Oat3�?,NZ"/�4˱\�Q��O�c,�ԟ��-�*���C0kX��*��Tަ�[�*":�zܓH��=�M��)m��-0�9�`�q�~Z��"���봓
qѽ=�;�-���Μ��&حLvaì560�o���By���whU;��ٸ8@R���|0�E��4;�:���#��̹�{��n�Ya����@��s���Q)	Z������7�'��]V�����;9��߸8�W�"�{::*,7�r|��ϩ��˹��=���ٖO���{:!˷���p����U��W�&庹<~,͏���+&�X 5O�s���).���ѝ~��_S�_:����ƃ�ƌY�t*V)s��{Ս���tC����=�(��cN�<���$��
;��Yçȗ��
��I��%�I�-���K3WT�R���B�6~nqɰL%Hw��;9��I8Q��<D�d�F�@�w��k���(ߐk����O<_�*�Y�Rȭ�"e �������Vפ��	����������ކ���"�����aح�y�o�B��x����2nށ4����W��%\#���8��3�,��N�TZ"�o�U������ͩ{�?�������-��+��_��~�=
���C�+�K�S`���ʌ�� E����(��k[;,�Xv��s~ƴ6k�>���};%�o����;�m�X��'���@`�O�$���LWO�h�F=6�.�H�5?4�+ �o}�4j�]����J�'Β�풱��
��5>\,.4�V-�Ԑ�a�H	�b@����V���]��݄�X�ʤ��tN/��i�)�A�I ����_Ԑ��:�&j"g������M�q^ �4�WG��"�%������u��/��`E"{��u�D�0#�'�@#k��f�}ӗEp9��ZgLtO����v?�PL�t��ﾴ��P�*�9�d�L�KSz��K<_�@չ��q�	eհG�:~����H)��7g�A����8��,���$rnb�^��I5�]����S���k��3$\^���7}�S�h�P�+�yt��Q�ϑ�����'4��q�IQ&ۓ��yk��؋��a��8�l�����<���nCK^J-UmD��y��7����\Y���߶]������^#�8r��*ƨ`Gw����Vw�+��-�Q}�?nmс[A�NteXu�6k�cT��`taMs2�*�t[�_�y^Zd��� ��`Yf_Le5<A��>��f��S�l
At��jF�`:�y��Ɖ�چ���r9�k�!�F�&N�U[��%�Lᄢz,zVu��G ��qd�	��� W���Z'�Q
Z���:f�h��gbs;;I3�����W��mA/Tot�J��ۨE�<�pߎj�\��	�!��q��ZuV�:d��^��{�i_K�����d!G�r��̀'��0��O�%���b���p��udJb2t�&���m�"8�"��zTú��ij�V�i*���s�n��NqG�t�n��aK�E�������������%6�/f�����;�á�z'�}fDd��?Asֈ���[s��: �r�t+is&RLx�(-�0u���RxX���g�o�͓y�TD�����Ň��: VX���үy�,媷`�xv@D���(a����5��sJ�S7X뚇l�>���r`��nm��%��j~��H���+��b�:���j;��f@? ���e�
�2ңxvy�Qj��딽Q`^��՛�� V�Ī_�$�e�H�ˊ&ԣ�-�N�\���>���uW�I-h��VJ�l���>A�|8��}X'�zD�J|� ^�>�����-�����Yݱcp���V�����>=9��w�'6	H��&̼��:5��Q`_���G�<�.�S|��X�Zaj�,�C&��1���C�c�2wW↶2`?������h�^&�<�`ׁW̌�7	�qK���V1�9�bt����h{T��o�	�p�u�@1��0��7����-Uep�AM��Pa����O�9F�1�Ba���$��cxBe���Q䰿��e*/9���?Ft)_��A}�n,yc����Y�/0�ukzi���ę=�R%�B�jˎvIgB���*e��d�ˢ�	/��]�M�j���d�����&���DBB:$t�&����2����h{�f�2�A�m�UH�	Y���;�����=�>�� 5��s�cYx���&ԈÌ��a5y���f����
���p��I-+lm��D����	ڸ�o118�;u�E�FA˕~��rw1m��h����A,5�(u��o�	Av�2�%�2��倐B����	��OA>+H��.|�i"�����<D���̨V���,� >��v}�'�<`��!�=R 5�!�T�H����.�g�r�`.��iw��x�u�ρ5��_��2_4f��j)^ry���:V�ؤ�������V=�4r���LJԒ�20��樧��<�~Da6)�m6�$`�S}\�5�r�s7p/~TS������ȃ��=�rr��a��mk�A�P$��2m��h�{d�KQv�ˍȡp3�fa�k��i�+92p���_���(lx��߯-6�5��Zd�*�t�K���Mb��۲�'��qB\r�5q�`r=�/���N���Fs��ݹN^.�bd�m�c��n�7��{쉳�17���vń<�����Wɮ���BZ�Wrg xH ����G>k�*ý��]5���Ɯ�ֲG��M*b\#���]���ߗ�T��
�W�J*CO_7<���dC��En�	p�nm&�����J)F]�K)}��=�P����#�AER��f��;=]����:�l٭s�Z�52t�t^L��?x�àv[������o11{SJ��^qz^0�M;v�(��dU��rO��u1�,��-���Qn���h�Ur��� �?E>���8�=td�@��S'�����$�$�f�*!��H;Z=\q����R�RxF3��h>�J��ܙ�l{�(�W���΢�fu]�6�^��,X��l�@�7��r����>q��x�39aT�� H��di�@v-����h��ʼ�յv���F���>�3b,r�pȉի�P�Z���F�lv�`��~v�wP�\ZK��3�#�Lٵ��K�ji)�^���|�2���#�!�s�Pu�C�����M��z���ŋŶR�yhY�p�>;�����1���,�}k+�M��LۜIn����f�������k���=��sa6h��̊3�D����y��%�[�P��Rb�8�c�"<���G}J�������upn7N��N�sR�Ie�j%�y�-6ʠU;xo�Ky�;����T%q4���8�Ҡ���ABVsL|<Cl�!Ƒ�)�X�e�Zw�;�wk���Y�#X�� �w�B[�ÃwY1��!���^��r�#�[�
r���!�A�������C@CU�����n<BA~���b�1���b��Pz:��CO��6��]�s���>�Y�«��S�A_�XǺ�G�}�C�������装���4���)��� �Pw��Su� 8ev��B�J�IA^�� �G��'8'U��-|�u�5or������� R��R�Ԋ���l��w�s��:��GEf�8?�uǹ��kka������ڃ�I�DW��Rk�|�ʓ�T�z�s��[�3ʍ{��:fB�������� d��_�R1[I��d,>1A/�&�<9�1��4��%x�K	]Ἂ�ȩ��(�lw���z5�n~S�nK���hq�O�b�ʀ9$C;�{�L��5���^N����q+R��&���x�n�-��Yz�Q�6�Z��&� ��+B�@��SQ3���(���ѹ�&{�^�&	�)�ۇ���a��,��*1N뛢�6��CT�/Ƣ�:1��jd�K\����S�o�@$/�u�������p<Ecv��$uTY)��r���g�)��V������WQ�G��8�L��~�Wu2r]����bv��B�0� �넍�ک'd�L_���.Meu���A��.���'����A�wTR��������}vrLF��	���li=�6ܶ�kw�C.��r�?nʫowA���QG߳�Z�6*{@{��V�c���&�l����Ld�P��`U��?ٰi��n�\�*�$��\��n�/�r�am߼��5-�nǨ�z��wR�;�k@Y�ޢ]���9x�z�T���]�����)��l[ɓ�g�m�-+eu峿��Bm��?A@EBU��3��i:8И���t���n��Jc�<�~F}���XFN��E��K�����TԶ,���NS3#A&n�E���r䊶�
!q��^ds
���4�,ۉ�	-�q���!kd���0�"%���7�q��I��������{"!韣`���R�Hw��Zk�A���$���L8UO�P���?f4̇\*����M�`�Dfֽ4�ڗr�9�5�C&���%��2���N`|�
l��{a���K���=�}�,��v�'�G�%r�4|��TDV�-�;�����`&�H�,�\�Z��F~́��p���ް[��!�h&/�Nx����.<=�7�`�0ƍ�}����zD��R�Y���:�֪���"�G���q�nu�����:KZ�u�M��V|.H�KU>�M@�`M1����~�.Ţ�rx]%���4gP�K�w���/�2�Z��g�>�:(��]�.F�ƣ�DWY���*£�6�t�|��ȴ�h�;��ǹ�d�MaR;.��lK��/��C��K���g��m�_���3U"B݂U>�]oW@��@���r[v*-�dt�3���� �����n��ZR�$�.c����lL	w�&*<v� �u���og�#3���M�κ�)eE�V���6���|!�l��{R�6�^��,'�j�����L�Yɻ*@ ���8h�n��NZ�|���;�?�������J��AS_�l�*��!`��,uΦEZ�Vy�"`���z^5�=K*44o`�o��Yb�K>����{mx��FX��� k�ܟ��41`n��v9;o{����K�E���|%UF�2,"@���V�)�������}�4�##�����"���rE�b������Ŧ^��;�:�i�߫�z�o�i���/vW�i�r����ɻ�M��F��vrرݻ�d���3o�!��T��m��>�ܿ�ibDfY���bQw4@HK��_���; Z_\������IP_ˉ�x>�P�ye�uӤ���YCdV�rf�;�$��ВRp�DL/��TnI��>�����@ED��IՖC���(�Q$�Q��<t��O������%r�F��%����4� ?IA$h���}
����L�QT��w�r��>��P�ϫ,-uV�d�	pg�&���.@���'�Y���8������������a3�(g��ף]a���ݍپ� J).{�ђ�"Ka���=}&�%Z6.�#|�+/C�t�V�7Z�:��s3(#H�������K�������fMo{���0.pY6S�^y�zG]�a@��-U����E���QMo`�m�8�n4i瑏+n��~
�ɝ[&�.��8��K/?���'���9bҸF���4դ�#&�d�&����̫b�iZi$,�z��*ժ��_h��C��,~�SHɾ�;�_�>	b�G�-��A�tS��6�4EY|a�����&�z-�	X��	H�LY<¿U�KFG����[Z���:x>1p�Քܧg 9���YMqy; �k��&�{xg8&�8���R�����h	�خ��@��P�T3�����{\�)V�Ք��Wq�s6q0��^bp�Z�@a;
7��y�/��dPez���N�ȬM��]|����ti���2Z�6<�~5\c��(B�|��#�B �ƒ�ԋ,�-��c�J�&�iR��C��lE_�*�a�yQ�E�3{��4~4��Y�����MHnʋi�6Bd�RC�E� �L�{+ъ��rb���[�ɘ4'���#�C��kVC�*�X�#�{�����Α���B����o�c�Z��#��]��T�k��q����{�4DlEx'�HU�a�(}6ן:���h�{:j"M|yR�m<�.��T�7�x�jG�םk�;Y���/����(��-� x�w��>/ 4^�yߗ������jB����1�����6�2 �J_�IXLj�SzE�Q�����p���e��`��`���#fPr�l�<�7�B��w9ԡT�8uE���
���yn��"�]��	�#�q�3
��D� ��Qb�`�0���WD�ɘy^�d�0?J�N����@��]Z4O������R����z�拷u�~�������s:�H������}W����3|jq�ځ���U�O�b��f[����0�;��xJ�(�8 #���7/#�w���P���'4�� ��V�F�	0��l���L���7a�YJ�W�x^k��*���ƛӺdILJ$`�2�g�ݸz�,頲�l? �>u�FL��d��ۀ�Y�.�����F���'�F},=UP)G�h����!B�o8ª��@n$e7�8��Wl�)���_4G���W,�+�o?���Ǔ��@�`�M�ۇ��Ť&�G�2%4[m�B�Nz��%�*��~!ք[��� 6�b���Ǚ奘������v��Fd0^�H�l��4m�±�cN������`O+������FHX�@9[.�>�$�W,fM";�����S�x7��_�i��'��(~/�D�y�bKz�wE�����պy]��	���çV���������N1����8]B��EP�G_P��{8&S+���1����jm: ��}kGDG�q�kN�����?�	피���)�%~���v��&iؤm�;��oIE9*_�� 38��D�h����U�P��K`L	��*���[��*8k Q�G��hw�aV��/+�2s
P�7r4h�;���s�t<�GA*���c�J@9�)���W����6ڭ�z ��XV����RoGJ���[(3R�h�]+���Q��v�Օ�<94ѿ���b%r��R��xT����(�N>�-��V�)����}�A�k ���ր��B�YH�����r1�����hG�3�=ELY[�@��q�iq��fЉ(�����$.kQ@=���}���q*��n�^i�Q����<���˸�
���j�C?�E�nf�X>�q�q����ZN��/�?��R�\��]�]	�u@�P)CxؙRm�Q�8.��
�|�W�h�;�ؽ�f�͇QU�Y`2�xJ 7���}��k$	��2)i����'[qAX&�ʍ5A�EywY�v$];~�ר���/���R+���;�e.�3�:A��?��D���m�N8�.����a�Zi�?H9)G��ӁH�,g���P�Mf��EA�
���܉>=��'�hE�ؼ1��Ntu�+c[��Y���˸GD�59`n�`h��[��m��[(�HL��8��_�5�gbj@�:���ؗ+��S Jp�Ǭ&m	����ŁK�p|or�G��7�O�?�OΛ��Nuz��.�/,T,�ygZ.7qM�R!���1#h�����Z���9��t�Q�Mm���z�#�<֌�H̴&�n
	��Ƣ��Z��r��-��Z�����O��!�7���~�� ||�,Ry�7_���6$�*��jjc_�>�	e6	A^4�Jq���l�4|�fb���A��xhMD�;�O�����|�fצet�W���h�]�;]������\�bQ���/i���9�h G�\=R�U�����z�� �_V	Ja�-1���o�/���;�)��٬�������#�e>��x�ɪ�AE����H9�d ����󴺆5��m�uM7Q5��|��U�ѿ�$]�2�Kb�B���W���������$�]@d�$vJ�-	�*������c<�����\
J���n��=��b˰Q<�(CQ�+�����Zl�)�����N�k�ld�UD��5j7����_�1��:h��4�}���
�,�u��-��W0��Y���Ƥ޲E0Vb��쎭:[���� 3�����ڽ
f��e��`��_����)���'��R��=�`���/���[8��)�b�&ch[٣=��l�@��h�ㆿ!�ZY���PFd\Y��8w�/H�E�Z<(饷ZF���o�J�S^9��.D~���s �N��6#{lj��j{�����S6����\�<1푳;:�ٲAU���$�����2z�g�����<œ�m��	��[��/ ���� ۘr9V9�M�:�("��[�FИ��[,.�^��
�S�y�;��:S�:�X��T���m�;�Sn�v���#uqA��-����4ɋ�,�������5�������x��f�Wo�w/����n�W�s�veP�����g#Mg,�9�^�yp��&M�E��軃 ��=���{�b&ܷ[_���;�p�� ��2���5;�t�/��>+��:�p]��1��$?��l�
 StE�C����� ��'�9�J��aNr���s���X���Z'��(�}%�[J�e����%f����X�����f@�b.�����F!����g3�*q���h_�qF9k�]c�c���Y�>�2V6چ�_�&�s�4<3:�)��3 ܢ59�"��b^8G*� ��7�F�[��h��ĝE���o�vo�f�0���_u�rU�)&q 㼇@��յ��N7@�e05�Y��8Ք(*{����)�ypK�Y������ƚ��@p}q��I-;匵Y�`�����L��.���>;Q�l(��G��3}a���՜ɡ�E�����ۧq�z-�Sh�����a�܆KT�1J��>D��)�8���%�s���_�n�CK=`N�J�I[M���jOtGE��G�úIV(�e�U�&o2%FԔ+P���>|RgaD6��)���?�A`�f>%w����r�LW�^r�&���k��e͹�}�R�<�~&U��M�<�9嫚o���L����M�����*����)o��v.א%���V�z@�#�r�%\}�{�����5.?T����?S������C�yښ�w)'��0~�����ބ�6I������L[����������������6;�E�l`?�,�q��Z�a��Mh�x��w����n�1�\���s`�J��+�~�l�l���1*�'J�vB�1���yRH��`�Ͷ���Uh;L���+�y`����n��3x"�G �2�
��AJHi
5L!�v9��ѿ��E�E��=��(��7&s_�h E9
Y'�M�:�Pd���RV�`�ytWm��؜�|��&�"g�'|}Ĭ���Z����jN��i;=��cV��sH��j�M�5
I����8�EAԶ8:*����n3�߈�L�� �"˽�M�3Xi7�< "w��L�{S��$�T>��"a�cp�u�E�r2M��uk����'sC�q�Q�� Fk�Le��8;�?m�e��P�*H'���5��'a�9�k��7y���$EWt���{޺��P�1BE?�%7(��x+�4ڗ�*�)��!{����`*	�F\�Y�=��]������9#F>�+����3A�������YU��i����\�A�??�%��;.��N�D���@zWq��!�c��`��@�s����_��,Or_D��~Zn4�F�v�GO�A�P�
F��.S,�6Հ>�,!(��>F?���������5Ξ�h(!�o�k~y���t&^9t��{�q0�/�q��,�X�o���p�=|��Je`�gw��;򂭂�����
:�Q�a�15jhqK򰡡#DN��])��?f�����
`�/��M2�g�o~ݨ�r���q��9<r3�>d��$�g��RW��^�q�m����a�� �l�	�
tK9|�Nk�0m֢_8d���~��x�Ȓt�VD�H~�&�"Y�_�Y�ћ$��V��t9�RA ��в¯���֊i-����6��pL���`����4�BD�<�Eu_�w��/&���:lk�x7@Z!d�S#$ރ�B�C�.�#đm�"�Tr��	HS��:WK���6�ןQd��f��w��K�[f��q��Z�jKY��a��T�x�~��?�G%l��$�$�y�@	�/��P()&ϱ9z�ĳ�V��Ng�1fo*�B@��զ�2�kI�)B�v���ܧC+BL�*�ksPxI�T����A������ͽ#�_�nSڐ���-���0�oy>���>Hښ��i]�H7�$F
�^�<E�_e��i�s��b�]1Y�X�����
�JO�2�,Q��9(m�H�i�/S��[��^��?�"�
�y
�>i��`&_��w9p;8�F�g�,�a�� ��
�b���M��bc��-��Q��FxH�أ��c\hz?��.8h:ƒf����a��x�3-%�^�'R�H��P�V�.�f����x�q�)�E�뗊G����~�(ѵ����0{�A(`4�S����$�N�����RЩŪ�]3?s��2�k���X��Qg��Y������'�7(��(ǒ��B_����kK�	IȞ�������a6��D�bW�w�������=�K����o>��Hb{P�M(�@(�3��KV��*mQ�GI����`a�M�z�V��.o �k��8 �MogN�!vx|p��!�G����C��B&j�&ߘ5Z�w��o)c�Q�<d������]c�.f[]���ߞ˝b:0N�4� ���x��b�Z�A~�D@Ms���֧�������qp����ˬ^��^�w3s�t��3G����%�1 �� w��0���6+��{�3&�]�l�?,��V�b�Ϸ�7�Ih��q<f�.�]�7W�n���n��h��L�G/�Q����^�r.��ngPN�����1ِ����aa�{�v�X��d��&�+~��6���^n�A�H���7����&m3?�	<��͕F��PB�_˭T���^�#���n+�09k��fH�� 4|-��}F0�	/9r�kשL�������ܺL7��NR��Q�]$�'s>�G��ǭ�o`t ѫ��9���]+�P8ā.l�����,x+�����E�g��������~V]X鹣�]�]�����Wj��e�g�kJЬQI�`��W��I4�_+�C�q����~�kF���Me�e�s=��ٵ�Jle���� E] �9�����-Z�����\�f�5þm�v��9�4p��z�*��1�a/}M^;`�%?8���O�Z�p-��t
�:�9b�t�#!~<�:V6t7#�L�"���r�9/%n/5-*�l�,AO��7!ʇ�J�ǅd�1� ���rA�+w�J	���SI��4��҃�[�U��d����W}�jj:��T�J�1���~�;�����?����%�����!�q�5���������c�`��?:�R V��{@HfG�C:A'*��rCW�$P��;8řA���q ���H9螖D<m�t�1���)�x1�9�ԵMM���.��9j���� Ȇ��&5��Qc���՟��
����1������I��Χ<���R�����~V�&~a��SZ��3���=<�K�e��l�r!?C��R_F`�f�JJ�FdB��V��9Xco�Hŀ�d��~�E�� �h	��(x����eD�L ����� %꧿EӉ}.�%х���_&�)!܍��z����w���y'2�� d�����6���xO4�#Y�ǡ��-�$M�;�����kg����o���8�+���c���0C�i>q\
�'�;�$˰z�(e-�0�Z�u���N�tk<�	����р���F���9�je��N�~�j�!�U�Q�*�@��$CפŽ�L@:6Bf�;02yܾ�rQW�=����]hɀa1%a"�L9�|?��0���/�כ?�`��XÂ����R27�<�Voi"�����L~�k5O���`A�X�͌���-rs�J,���-FD<��+3�3Q0�'�7h���.h:<���&l˳��&��D���~[�<�f��)t��6m[ᓖf$������h����Р��ZКj呻���a>���p�,�j���Q���t�������<l�����W�:�Eq3+R�{<�����1�K�s�ԛ|L�/���<,��a_3 �J�Nz�8���Ā���`�U�K��x6�1��KBp[�<.C�&�9��L��G�y?|���h(o��g�c~a΁�XV)b�4�5�EozX�{��8��`3	���K1��
��a�y���A1���5H�@WY���몽���u��+�P^�hq�3�O=a����� ".�����aI�+��M�=����cu���� A���G�<AG��ց7�����B
���4�4Z�f�~�f�N�t���ƚ1"$zEp��UD��l����Ò�����b�w�ѫ�L]@�d�p�xĜ7q̳��'�~��ԍ����a���L�{҄/Z.D�l�ʥ��q
�+3��K��k�[=�a����W%�`݈�������3ZFӺ}���
̉�|����s�VT��=�)��Z,%�Ԣ�Ҏ�`��v]O��5����6/���@GA ��>駸����-����c����9�d�`���m�ǖ|�re1mU6BԽղ�x���ܫ��3��Sm:�c�,���"x�J�g
���dk\c4I����Q�Zr�$��L�Lp�/�H_�z����q��[hm��w�0}�:ܣ�t��3��e�/cs@��%+�"�V�02'>��ǭ-�]�o7����l:�4d��M���̀fq9���D��z���?�&��*Y��(׃�"���|�4=k!�e͈ћ?�wI�{ɝrK��.(!�洙%������Z��9l�tr.�}��������fן���@��k�*<�@*a�������hnZ���k�b�F�MK2S��?�e����.3�G�o�
�V�:=���#g|���U��v����)�9�|�Z?�,�9��I'�y�Cu�:�S���ǀ���4�N���j"����>�	x�3c`�� ��I71Xx�p�� �m�G}�+|�m��-�� �I��Z� %�~��o����0����������h�~mȘT��Z'(NE���vW��9��m����E95��Rm��'5K��`��ef�:w,�� $ 7����
�ܤM��ܖ�g�1:(%Yҿ��`��C��e� �u&J�W��8[@L�!"7AY,�;$�s�[*�Z(�+��� ��/o�b����W�ӓ�|�s��u�ޘDH.0=JU�������QehCs�x�ڜ���Wc��5��y����zH�v0�
vX�mCP�J�N�#=�C���k?x��RV0�yj�eF�#V��FA�e9����{������R(�L������q�T�g���e	��������\G4i���h1��nǵ���FM�\��}���,���k�D���b�Dw��g/���M�@U�΢�y���ZJ��gM9�Nރ�������YB{�q��K�l�ԝ����T�`!�����7}�6�12$�w�)����D�|���g�JrN�cAq~ݪ��ګ!�>����M<��^�L1�Z�SKy^�����ܛ�V�9¢���z����Y��,,]TQ���� ��k:x�E������8o�/�_�x�m"�o10�T�=s)��?�<	���2�O0�1����:����<9!:�=ص����M�q� |+zt�Uu��a<��,��|)O����)���G�lŬ/�p�M���}6�����T�g� a�X.t%�5Z~��e��C˜hS,���[�a�~e�X��i�A�����m���:�X�xMq�@׳���=$��hד����W���K�G'J��hp�MI7�{w�x�݂�שE�g�M��{���	�wk�
(x��Pi���������a3��m������':�<e(�(�s�X���o���1�����)%�d��A�F��Y�6=�OY5c�靺2=���+]��j9w�@�4�` �M,��n�F�S��Ǖ����a7-x%8I`i���^��Δe�q"�!ķ�Ɛw�� l'��fR��#�?@ުHe0hˢ�����h�g �5[��8j~SV����@���*GY1~$�A��a��q��b#�H�J����@�ܴ��������PhvЍh2�[t�ͥ�.��K?e�%���Um�~��߄g,|qHBs0��/}����i�k2Z�~ ��6t�u���
b'�2��#�ڐBgK-�@�Z�gH%�n���S#��ܿ��o%jei�R�|��	� �p,1��o�cl�b���}�d�ɼ�[�Cm)�ˋ̦�u+#tD~�.B
q���&]_yo�uNϫ���p��2���m@�ce��M�]?RP@1��`����IQ���I&:�9�"KF��	���>����;XF6�x������tg��F�GA��S���c�����m���Ɨ�*	��?2����W$ 
'�W+��2���^��)us����KY4T"�Ҩ���P���b[���F���ޛs:܊#��m:���v���/ky�n���|v��5l�ۗKtk�w�T��a�R3�Ts@b'@���>�J���ܚ .�_N=�A�k�<H����=�#C��!�"^��ސ��w-�HM	}���n+춤���ND�u��0������	g��o9nލA���,���AF�͝�@���xb����}c��O�a����W��G��T���&Mb7��IT ��p�Q��:trޛ�g��k��s�]ס
�he��IG(P:�5R db��1	$�8h�x�7S��J�Dc�+�UH��z� 0����;k׆v�m�8W�@�FXڡ�S#�;O��Xy߰=�Cܙ`�X�O��`�%���w�x�9<�(A�P�!�I���պǜ��A���;�"�_�V�VՍ^ �����m94�b��d=�+��2�5���N�լY<�V�y�{����9�E���1=⁮�@s��8�ٍ�Z�&�je'�m��a�8�%�o��\�����������8�d�p��WqӤZ���`*:��;����m�Q�0U��ۖ5�l��0���������M�+�{�)4g�
D��˧JB�@���������IE�(�;l-����.@ ,�A�x��BA��;ݢ3%���ٹW��~�t�i����xU����ᯭd�e�.���I��H������4�.Z"~����gX�}{v�)F��!;荌��H^S͸����*ۆ�>8\�tfG�{{��ٛm{p����]Jq�ZG�|��.{�)p�l��$]Jv�;Í��c�4`�e?_�ދ�����õ&�wLL!k����咓m*q���ٔ,�FZ7I3	��m��q?�);��0�F�(�܍��!����CW�Kv������C;^Mˣ����*�um��CIԒ���G����N9�i��2�|�>"�qt�U~l�sH���Fy��x�4_�IC4�׬��S��Xm֘�9���<��^;����ܑ9������z�|M�P���V�@C�3�ܷEyл{��7Y����,B.(T4Q�Jdt���h�)�s(��}�M����xm�M�%�)I&X��ſ��_x1�On�T	d/Y��޼UXbK�v�Y�[�V�@�)� ��.Wh뱸^�5�$R��?EZ�Tj��9dV�<I���9y뾳�;h]�5��P�|��zC���/_�����D�����nF\�f��9;c��^��t���\�����m/��Y�T UX��w�@��W<($*9�x�� vL�M�f��/�1�u���Q���Yй��R;���������F��j���D��/;�ھ���Sc���/��PAAa���BT���@��I,]�*K��몿��+�(�D�^���[>�\_#�Z�
�Y|��9�GvS;f��oq���"R���fk�@�І�K�����g���5�'aR��홾bٲ�-��zS87LV�(L�V���)�א�S}�U��σR&�8�u�9��e��	ŷb�Q�/dXY+��[�&�l<,�����ڰT��Q}W�"ғB-��m�[x˕d�:eZ�f������_7VH@2�Z��>n�&ހr~H�C �Y���]��G����e}�]�[ʽ�l������%�>����k���cS�U�U0��np{��+���J�S�j�^�]r�I��/��NU��bj�s.����W�;�-!��]P�3\'� �g*y@%(U��sb�c�;#�J���z��u�i����t�-�'j��\I?n��"βL@�I�Ї���A���qR�����|��6V��Z?V\���T?*�|o<���oy�[�Z���ّ�,2uŷ#p��)RO>A2���;����&������$��#�M"j0�˾m�e���
�b�o�C�����f�Y;Z���i�e�����1�ڐh��<�TWݤe;�D6|�"+ 5|���k'��L�q�&�
��	��k?u�{=.o���	��I��7���bT8��~U��'��n�Q��ӎ_m&�E�i�١���'S��<�P�E�p�=���z���Ɛ$�}]5�QvB �O&tc�.S*�D��@T<������wW1H�O��2�"�.�xh!�X�<�HoLǽ�v�1�_��`�(�S���1W���%�%�Q����$���P)��Rɽ9���4����W�U�9�X��dmᴖi1�	Ƣ}�R�/�n*�$�7�ӆ�o�.�~9�*#8="�(��
D�򄱧���j�48�ayj����(���hDg��W��rǜ��n��qү}
bK,��)����"j���*�
\R��e�{�H��C��y�C�e��.�d�v�>�� �<���]�g_)�)�ĄT)��W�6=R<7ƭ7�!C�gyK~1f�^_/w����
��G(e�ur�O8�
�f� N(�����8�ا��dd��Ks���C� ��j�倍1k�������<27����ߒ�8�+��-��w0�\�s-��èٓ�X��.5�(��� i���`<�cG��R�YJ���9d�ji,6��thŉ�7�m��� �CX��q3�BO�2�ؓu�l�� B�eM;�PB��L�dAa7����Gt20Yڥ	��%�)���m���D�N��$.@��.Jʲp�vȯ7r�ccy����	w���ڥw����+8����b�h���2�a���b��"c�ܳ5I���J��Fo��Ƙ5�<"�9n���^^Η"Gt$[g/��4=79�[�S���Q�'"E�+݃��Ʊ��w��k�f�ܲ�_:�[#��s��2a��\l��ŻyF��T���Q|��T� �:�z�lI��ē�.?���#��(r�$�CL����,�6`=j����ad��"N��ˡ�늃㺛��������.[��x��Q� |/p��|FOy
<���laZ6�k՗nJR�>��')1d�������u���7�K�'sP�Q��?&y"����{���c;5g)�C*��vE�vI�*�]ƈ����ݝ��<�giL��L��1���s%P���e{�.SY�)�1�A��i�$��O�������{���nCk]��"
���$�V��'*\8�jv�	�Cz_�O��'b̀ϡ�[�e�VW���[˯��lP����*�ڴq�zx��O7�'���;>����1%wz{+�,���w�]�D��G	�@R[cj?B0�k�qau����G��m�3ڥ�KX�N�B,��t�ɾ�0G��??�#~b���Q�-��̃D����#8@�yoq!�M����W��_��D؂�Б`C7}��Gj�2�Ɂ��)���=&�^u�tA2jzӳ��c^��8��-��gS����x��I/XƞF�[��K������e }����#���<L@.���=�}�����
p��:�2�u~$V>!��0����:}��u��T`W}�w���g�rwj.ڳHw��:��kc�ޓ:m�~+�s��m�S�6�#}�p{�V�:���E��Oc�R<۪�|){wb4)�A�n���k&�An�}��"6U�x;����M����?������! �f�W哱x�|�+�~�Ow2�
�RUz�.�B��(y��▚�`8g�iTh�Juǐy4f��yc�|�#�_sL��6��=�Q6I����H�7���W�H��w�q2]�p�h'�ei�ec��$銐�^P���x�M�W�e��%z֚�%G�O�X,^�X�U��&�c�/���Z��8�G��A�(����8(x+Ý�Кg����ZJ���s-)�:g@�#�5<a;B�cg{��漋Yo�'
p�s�KQ3�����Hk�g��BVֲ���*Uթ\j��J�Z��\�'-�ۭ�]�а�*9�?���g]���ƧA�,����ojfLl������ʣ�T�5)-�R��J��z�Xan���d��!�C�]�*JRܤ��fG�9��;DمE����``a�)����x�Ɯ���Y�(?�ɾ�����H���O  �<ݶ�(ac�Pv{d��~=�c1o�Tr0�o9:����lBD��0E��A+��u̓\���3o�k~[���Wv�YV!B�\�d$N7�d��ZVK��⼰L̚c���#m]�A�����Yd��{�+���}���F�J<���wX*��:`�hW�-(�h�/ۧ$o�h$緎D~��t40���K�3�k	)��o$OBE�%��Hw��Udb(Gɾx��w�aR+�!� 3?�J(���ݚ��i�}`	�Z�*�UI�z1p��¢���q��5ֽ{U9c,����^��^�6.�ړ>��e-�B� �/EƶE�"c�g�s ���w��p���߈Н���4ʯ!ʣ���djWF�}�h��������o�dn�j�0�},��Ԫ���x{�#I�C��������0�YG~�g�9-�%|�O�����f�v��1-�fb�f��Λ�q�Q�NO�۷�S�Nų^��1'�c�g�s�X�,��Π�lC��;Ў��f/��ǔ%t��}�?09k�}�M/`�%8�������X2	��"*G_�<�j9!�P*�I�oG1���9l�����IP���ʚ���(��j�Z$>��1���fq�AW��AR�B<��FP�������M������R����6�Z��;�]� �������m��?T����C����Ә��ݔ���B�i�5V�}��L�kX��0���),�j~�D����>[�;�� ��W��璑"[�Y�	)��36"=�	 ~�Q����� �"���f��Α�	���X���ܤؔ�i�_��nh�e�ޢ�Ԋ2�<��4�*��Q�� ��C~�{��^m?>��R�`�Kg����nOU�BB#7�j���DǬ��l�s��IU@�i��?����� ΘO�<e���P��Q�Ԍ$�<JҚZ�h���q�a����8(�	�]]��T|���u�_?r5tד�5�=\��Zލhƻ�Ӯ��f��?黐����k? ��2�H;���%�C��N9�r�	�Hol�g4�w^�@���6���>6�ƕ�^X1OjI����8��U\[�&z��i�7��4M����Bw�T����֓���`L:�Np(�I�B��\`S�UY@��������Q�j�: `�ms'hyJ���k1_^d_?qEp`�	9|�P�^Y��O��/?��U��(5C�q��W�Q�}j�ڽ�S�Wh<M��6\�"��P!���/�ɺ��,�z�.Q���A����r���-̠W�8~%�C�?(��-�,����,�&Y'/_�k6��S+��hQU�w�Iy��d3����7a�d�a�wh����׳�u�r��檈�T*���ՠ�U�)�ۦ��,�gf�T�\n��]I�-�ڱg����~/�<5L<�	�	����91ddp �� �-dp��G���N���JI�J���o��e��-���:u��g��z��@'�f�w�����WR1&i���'���q	O��>;��32mqW�n��ԧ&QmG���y��Fɧ�y�)T�ڍ� ��il[��AU�.{]1X�1jW�s%j����P
�E8e��;�RN�5h
��(�ێC��B�=�A9���a��)�E�������"D_��/�p�|۽!-!,|a���p��� T��l��<�D�N��{|��l��S��k�����A�ÒDPֿ�v�)�%|��U��	��S�f��O��P.�Bz� {t�7`���$\;ٯ�����/T�l_����h����k���RT'�w�ʛ����M�d�g:	I�IR25=������ B'x���S�{��т�c��h���Љg���Pcɾ��u�7�q#_(,'�
��م����TN=��Ꮅq�(�� �;�"R��EÐ��J &�UZ�t��1��Tk��э|����"�wg�{���S�N��6|� �*������%�n��ַL�w������kH�Ǖ{Z �A<w?��jE_�w+��H�{���W�%[)�y�yy
�SMZ7Ř;�Kף$Xm2o9��B���)&�S�Ot��0{����B�D�W�3�M��A�5v�-��p�Eb|W�X���(�TڪR�{��F�>�<�x^3�e����6��bs��<w3����f;��vT�B���.�m,��h��zj�
N0���VFf�(�q ij����G@˘�Aӊ� %-\���2p�l�P�Y�UR���]`��\�0kL_�_�m��8�;�셳 ;kԓѐ W��D��d���p˕ ��-����αw0��ᛳ� f�x��
�g�	
��	�e*���)Y4��x�Do��\X��Ο�O�O<�.a�e�b��ԓmI�eõ���'����FW��S�ac#)��o\��8'\�w��.��UX�͍l��^<&�k?�L=`l��S5�߲�K���uK(P�a��"�G��� ^�+�{����7�6��2�lzϷX�~��TѨ�~�D��,�sU�U����	Qwj�P,V��+d��Y/��Ά��� �,�(��I�Y�+^��+�nj(i�]�/���:��q��jECO7���?X�֠Ї�eK� ?�^W�W�ؤ���5����ʠ'u8���C�~�j��[�E���46���5��cgլtCLD��ɯ\բ�¯�
:瘵ք�������9�]t�` �����q��$F�I���E蚓��f�?��*Y��_��������>ֶ�{?xV��AT! �d�^T��h�'w.�%sL++��q����*��>l/V#�89j���Q3.��0d�0�-I�6E���r���≿_���!�R�� �q�G̊�M^¸.ưgmT�e�����>_'�i߷n�����Nn:��	��@�-�[�z/�rS~�ޫ�΂�(D��$H\��g�w��T3�f+]w��2����DPORO!Fz��`�!S~ŗX��h���{2�� ���x��B}�<���_�e������0=����>~�'z�ە�$M��4��2�3�pg%����nn-�j=�P�Ӹ��C�"f��+�iه����Y;�Ŋb��E_K���[n���~�#"�)4]c����J@��I��>�qD9&:�v�o����:�o�	'xU�N�2��>���Kpլ-s;|˱����fqۭj&V�ׇ����
�vz�"V���B���e�1,�E�e�Q9������۱Ϭ�,Q��I���"8T��n�}�K�����$����u�������𾚂]6�n�'��k��ua�5�C��g��)װ��\H��b���{SLQ�&�(�������N9׀9��<�|4��{�
Q/=D���U07���"�t��+._zF��o�l�;ο��#�e��[bU�*���:��UjH��gՃ&&��5��\L���m�$M*�>w,������F�W  &O��i�~� L;����C�I3�b�D��;�}�꿠	g��b�(��}�n"�lXSn�L%��5�s)ے��hN�u��`S	QV��l{ƴ���Ȁ�S�} Y)&al�K��ѻh8w����=�	f��a��ώ���p(�L-��S~��h?�.��!XwRj;���wF[��;/b?���H(��ς�gJ�����X��/t�Gn0�'`�մwW)��Vλ�jwEd�x���4�i�&7�VW�Y���-1��_"������܂D�Q>��Q P�V��b�e:�X\�-�'�tv��W��ri��u�B��1A�B$����P�1Xa�=	��]�������5�ES�Zy*�{Ø���f�,w�_P
#O��h=W�$��~ng�����vEP�홈�O�mZ�_��ņ���%��u��2t�`o����_�M��f�fG��<����B�Ⱥ�l��D�a��*��7{Y�0�9�m�d����\��/�G�U[Q�y�rE3�����2CX�5x-ܘ�@MUS�ڰ���}W!�A��5v����1/wӼ�hv1�5N�U9��J�w�20鰂�'����?��\Rw*�FI�:,�	�{	{���Z[!�xo�/���o���e�����vX/��#�ۣ��@�c�kB�:X�3~s�h3&}CΘ.FExia׃AK��i�q �s�yX[�S�l�:<�����|Q�26�L<��N�9êZ�'|U�bl@=Z;�os�{2��ȺAh���y��СR4۱��^��t2��m<M�_���j�?������֛AF������Q�<OÑQ����ߨ�l#��Vε�.3Y�Z�/n
�z{��3>�	
��5���A�M�:ҽ�������4��)ס�΍R<�R���d��i��
=1g�C�cC�4�'�:+l�?TP�~,	��.�!�R�W+hR��^��@f��<g&)-�sﷴT޶s�E�G�MV�ڃcRq(6�>cR$�f���GD�9����i����Ԃ�t�S��{ˠ���"�EI{L�Y#�����<	���Qx��h��3�W����淮�t�t�
�E��9a5&�׸�Z��yWT�b�6�=ѣ[�w���K�~#��jXg��;�g� ���JC7�+��[��j���J!ѱbLf.�\=�/;x�c�����`�#���{M�&[W.H�J�ǐUI���$�M&�`�k�g��
8TY��0[}Dw7G�����s���'o<�~N�`�lYʫK�W�����;�W��&������{V�0\�=.JI�M�_�ċI{̝`���^OK�����k��pd��@��h��S�x�hC�3�ʹĹ�KM��",ř�o��6�w�)�6S��N��]�WQ ��I
�Q �0�6=۱/����N��$5���EQ!kBT!��o��b��)��f/fϦ�+z��*|��(�.Q����JS�Y��z���r��
aq��aqG�p<0a�II��s���q�i����x���Hr�k�TBL�Z����d�\)�r�<�v�F���x�\<�i�s��azsܡy�XsN'�8 �{V���;���3���U����F�j�e�h�����{c�aF�8�f���)�v�M������d�\������q=V�(� ���pQ"ٶq(���R$�P������Y���9�}��c��"qg�QQ�X]8<�������E%�HB��Di��=yG�Kv J�J���ڈ�5~�s�F�V]�R��M<
<SCj`�{���%Ɓ/aG���ʅLh�f���O��"��<�^�8wfH8b�����L9�5(��{nM���ݛ^W��I�u�^EO6>�T�T9��jqJ����X��	I�i|��7���J/�$dygr �.�9���sJf\�|�	*a6�P�_jB��!@l�A䰯0�ChBU΁�Mw�E�yWr�Cw���*�G���iٚF݃�5��y����5�8�g7	W)�l��J���FM��x}�D3DNS{T�C�A����W,H	}��$١�S-�]�XA�^��~��wq��v ظ���=���y3} �}�	Y�D6��4��/�/d�'+�^����4ۭ��|�%���Cy07{-�� �8]!#&̄��{{b�k4�p�S�2��۫����nI2�M��u�΋�+	�]R�H��\�I-���O�:��\�z)t6�EZ������KW YJ r#߰$,�W\�ތT�P]�4+Q.�<1M��(�<	
�G��3x�v�U�.]�ƹ���yz_�샐'w}�v��fɄO�4�^�,�/�f����Q�k't�j8.��rd�Q�b�]o�L�M�Bq;^�c)��P�&%f�0=���V�V�e֑ae�%�.⹮2���ۂ�����B�70��_#�cLr9:
�<?�?�uK�<��?�,kLrr�R�����Y>�y����֐t���gM�Rd@���7�L��7#_�5�����@��d4w4B�ӅL����eCA��
�s_�:�ȩBS)���f�2#�G�K�f��?��9�B�)���y}K�j0����K��i]Eb.)�K�7�n��B�2�5�����AWk�h�/t`���-K�I5�z"'Bu6f�W$a�S!*�*9�	|.u��Sّ�-�ݸ	����4M�a�5��6*Ŷp��-�j�I̀����FƄ�,��ZS����lc�
TT�@ɉ���R\wRN���\$���ܺ��5YŪ���r�93���Cڰ71{�����������t�5��"W����p�" �.q�ת���ƼO�?��g}����Z����(AxaeL���=��r:?�~���gvh���wk�K��8�D�;f�U�՟n�'}��
9� �?'i�}�Ű��U���"eI|��+��ũ���c�h,R�Q���ǈl�.�x��8,��ׇS�*�x��
�I����,/���؅9t�z��@�'z��䙝L��׽��q%��"�!6Q�,�'ܬWD�ZW�j�"��R��ddS��_OJ+�S�����/
3�!�+��&�{~���F�ax4m��6}	OPS1�q.�~�T��:�dɠ��t�b������[�l?�:��7����,�Z�A�	�zMT�-�׫��O�Ԉ���T㼍�&�!��&��f|���S�~Wb�$㼞�s\���v��	#p�q�g ��('Hx=��;O�"�Dq�2IC��P���y`:1��	�j�Eu�,G;
�M�O.���><��vQH�=��>�~���yW��:�M1�jx�t��-��5�<����fG���P�׫�r��#�+D�mq�8�M���g�MD� aTRY�+>0�x�5E%QV�.�x�{0�B�\D���hkZ�꺙��[�jaT"t�� QG}�����������y��*H��xW�Ir��Z˼#-�Dn~�`ݍ��en� �־�,P힭�.r[�)���_B{XR�����n��(ؗJ��A�Fg!(vĲ�K[��	#o�𮃲�EW(�ۦG����� ��:߆�TR��Zp*-�`c�q��~|;����&||�[S�,�)c���v�U$Da�?''Gy�:X��ל��Ffc��Tq pS�b=\�A��b�a�T�ߖ��~g祰^�7ͣ�͗M�D1x=��a�TfS���Me2�&�]� �k�f�O�D�yX�A+u'����i:�	�,���˷����rf���I.�Y�5���
.jV�tax�����z�<:�b|�"$'~A-xѕ3�l�3@+�`)6K��%�i3u�*�ř��e#��7uh�g �����<�◫�V,L��X�;rEs��Q�p���@��x���O���`!�f�y�Ɔ;��~���d�B��,�4�!6&�t�e�܇��l�"��-�S��J���0ɓ$����?�8�(`���g��G{{\3LE����6U�C�%Z�����(ҫo�Pu��v���7T0�&�~y�iʁ`{�~`4
%~�l�!&��J�+p2*$��YO�j����Pj�e��w<��+Ŗ���L��*\�����I�t�\���3����o +/nphq&?��?c�6��� #����_0#�&�d�T�p_ln��������`�o.Z �Td�=GgK&�fÀ����X�
qDxV����y�c�!��$EE/���MeP����~�yd��-2�5�[�N�@����6h.N.Hz޴ۏX}�+�3|��e�ʹJ|x7Xb���)�Ȱ��W~�MuF��㤥�4������u1]�E�*�Ϗ�b��X�ԈuVBX�_��:�Kr��x�bʻ�� A;����\�6��؁
w�/EŽ�w&����h��F�1��D��1W�K��^2�����͐7l�dr�4f�U�3��E��ZM�6y�+|q �,X'������LNq!��j�c:��Q_����ny&yOk�L�g��Z����u8@x.�M��M3 ���gL�1⁰�f��n�a�/�������\�>l~��*��t=%�ET`�B�lo�0{����~LOG�eH���1�M�H�}K�*�`݉��ۿ���at���Ç�l*9_�������b'�B������X���s�����/����sh�[��^����>	M�Q�$l����O%����~(�q�dN%M�
���޽3B A�^���([tSf��9}=��x3_GMΎ��*:nBe���V�� ���s�ϗ�����Es��R�#�x8��9_K�mX����|�d�bj�N��o
���)���u1ǝ+P�ą���X& L�U�R��o����D�	��^��'�|X�@c�*L�
�(�b��?O@�j8���_�vd�����L&�~���m��Ix.�R/�51%�>��2���t��ɫ��݁U��@�>���^�(}!��39�4���;S�Q<��K�dI&G������%�P5��
�8�\%sE�!����V8N�>~�� ���#�1��@��m/�s.��骚�(���,*՛�Q��+��oXK�u��.����0�Y��� J���J���P|LK	���o��H��=�+�^���`����6�ON��{\�2vV���ė���{�>1����R�6鰐/x4��(�x�ǎ����ʔ&S��Ns�)�yџI��~�=������S���?��I�h�۫�^�E����]W���$�ʊ��F�ޞ �0�1��t���<>H(nv6Ι��?/�AWz�A�d�m2�Y�����b�ǈ,<��H;T��� z�_����6T#��e���ռ�t;˲X�=�����0�Ji��m���+����m�4��*x������WzQBZI���$r72�а��%�E�QďE���Ojpe��9��ݐ\��x��%e�q��%~0���y�d�@L�zL��30� M�4��%`�w���UݮݘN]��U������y"��w��*\ȼ�/ɒr�@�DD4A��������|��ަ��q6sr�Gg���� ����$����xJ�����%�n���q�Le�A�t�_rr��(�h�-x���� �"ԒC�^�\�N�Y[���o!��b��l���*���<�a#��㎖ ��$V�U~���2PP�U��Ԯ����$c_k9��+���y��@r)m{����a�dZ}�+'xGv���WS[Z���eՁIe6,bA��b�Y���m�F�O�4	Z�0&�����F���E�O������rUR]m���D/JD�B���� Q�S�K��~X��@�	˲�&3�|�G���TŒHI�P�h%�ʛB������0:���_g����aЬ>�{M������f�����6v�in�{$��eƟ5n���ũ�`�G=�d�������@��ܫ*0\ӫ��.-2Mj��> RM��K/�<goK`-{����`W1�ka�p���$� ^D�ܺ�}v��&@I��$�����v�-���S����s4M�fd,|�$�{kG#��� �֔���7�ݣ=}��5~;�i�C釢���@ٳ���]�����k9����72�r]dYu�-_�V��Մּe�INTuyK����G�)y�}8�To��ڡp��A|O��1|�|j�]�����ԖՍk�yR��g�c�rp�p�l�s�V�δG�L	qW�$�D,W�o2u�M[)��a���|3��e���|��a���.��n�-ܳS��
%Y`��ĺѝP��߼����&^ĭ�S�afy�����[�nH��7�����=���:���v��i��3M|��7����$`wb!�7}k��Q�N�m�V�i�������8���&��0=�A�����豤�������D�;�����4 ��%̟���B��.�VY7��Dd�0n&�޽�]��3��>Ֆ8� �����7&���e��Ƹ�������s#���m��!7:����&��æ�Y�)��	����6� ���m8�+�=b��5� �+�y���Z?N����3~���`�������LB��T�M~C8�a��_(a��B}a'�*9l���+���L�Y]C��ΐ;hʢZ��*��)�28�=�m�C`o �Ͷ��n�NZ�_�zN��qc_JrB�촗<�Hj`�������h�l6��<��� �]���N�:�'�@�_W�"�畕8�c�J5w�,-ݝR�PU���I��y��쫞�r��W��:9�V���$��O�z�Q+6г�53�ZI���3c����"���
񓏂�gII��H:ׅ�u�B��d�!9/����E����F� �S<���N&N�ͪ�w��"��-�ڈEK�v�f�+y�C��#��q�,�F�v�?��ڼ�-y-��y�X �<
u�Z�EL�����H����
Ȟ\��t��� 2�~��	�f�T<���B24��eLC �!<�.���4��E����Ө��Om��������;�&�����ȶ},͔		u<)�a�	�Fи�H�0�D����eվ]{@K:�`�N�9t��e)*��|���O��ίgG��Y�9�E�!SD���&ȡ� �Մ^P�%��hLϐ#'�ʢl��ݺR�b����;�3�ͩ���
�,�I��Ha�!�:,bĊ@���U���O���k�;���F�>��|�=&{�$Lo�D"�(ҳz��:�4�'�>Ȝ�h^��+�dvK�muw�ȹ��[�!=��xUt7�/�U�]��*�l�Ѧ�#���P�7y��^�7FA�{C�dΰq�-�ɷ1+@w���x��:��Iۆ~ߖo@~$'L!��'�Le��{�֟��}����{��΀'Zߦ|O�X��4LY�-��Z��?�S�nވ0MS����.�-N���H��D:álUۺA7Q*"�?Xa@��,l��pi�I�]b����ڍ
Sw��V�?��0�b,҈ꓽ�����
N迿A!�x����60�ld#�9����D���M7����G��h � �G��m��+Z��b��(�4�	G`^�jlgǸ����ɋ�G��,y
�6n�~bEO�a���y갶}4�\�|��C�rG]���_��nTF80����K=��ـ�S�ۣGumJ-^1܏�������\?���g�vH7yY�2Ud�W��/Dd���?�u�iy�B��N;��S8�C��Bc�D���{�����^`��D����δ�!�'��5�$��2j�㉇��3����ֿ�Vc���ta8!H�v�!�\?rZ��"7�|9�
)Q��FE�q��k)l*�2����f�ш��7�I �"��r�f��%m�/*��n���3��9�g�i�w�L\.sE�!A�5�~*]���c�{K�Κ�A*C� �>��'�}�5�M�#I�Y��e�U�uθ��ɹ�)�?�����Q���qpoN7�(iX�5	�ty�?4�Q�|¸5��Wz�,C�Q��:�%-�k	�ohj[��W�2��� �{�'�$'�� 	�,�]��H:��H�ie��ErL�9���%�5w�Ṕ
��݃;�x�p�7��IWu�*������/C(Ӊ�q�L��$�ajO��f�u�&� PK���!�y0��C�v^N�jx�g��;�5���Ou ~>�l��z�K�������F]�b *�s�����h��O9SF�����7xH�R
�
Ow@�2�~��}���Дh-	�T��ͷ�ppiQV��y��kCq,�σR�͛3��
��u�an��Gˍ���"oK�k�\Q (3~�/�Qw��ɔ�:�};�����۾'w���YdL�b�M*����sz�*b�n<^{��
z�P��W'�r���m�(_G�|�o�a:�!P�	�a�߉xD*G���X�͙������]y.��>���!�t��z�o����T߫����w��&��f�>���� g�,��}s�|�u{i������ ��-K�%�o�}Z����n�M��"��NU�Ih���	^�9���Kˬ'
�Mt"rd��Q��+��,�)YainT6tR��3�����2��E��&�+&"�e�YTg�Xnxw�IM8��=�޼�5ʯs��(~%f�FR-�C`w��Ӥ�|6�>B�?|n��!��w+�[8��KB�c�a����Pe�'D�(�B�9�"��R���-+#�d�2��K��Mё�8.n� �V@�%� b@�C�;�k:���`߃�D�6@�p������R��=e�ك���R�ʩQq�>�J�A<��)�1;b�]F�s	�{M�X*\/0㥳�=E[��p(7���(��W͉|m:��IӗLK��%�#[ڎt�q�v����e�r�H����ti�M)Ѭ.Ϡݢ5���d�����.#��2�2Y}�I�1��-��B݆�j91�;AR��M쾲�S�1EU^�9�l��+����	���r/���v|×�8�xr����L��o�ɦe��;f8��c.4�}#P��r��jn&/Ι�4�L�9 �moK0qm�T֝,4�F��c`�7�a�f����b�,�%���#"� �V���;,}[��a)�>*Fj��Q	-t��`���[J?+��x�2�a�w���;�f����C'�����Fvݹ��JFF�n�i�PGPF���j$�fdC������X<+�P�G���h�A��Ш]
Kd�<���
12F�^�|V\�j0Ůy�^��W�9y�����'/�Yf�.��v^����5Ĵ��g��f��{��UAr�`߮�$ըN�77ɮ������dn�Ew��,�I���s8�C��7;?Up,�S�d_ď
��i}y�;-�b���N9�=f�i� ֦λ�"��N^p�|�-�.�po>@�L.�$�E�Q�b�C6b=�g�zf�8��S�����K��.:��.���~lu���&�@z{h���� ���?s^�#�mZٽ���X����<���3��CpBs�sz���d�F�(8�����.4���d�����rQ.!K�^d�8��޾?�!#�/��T����R��� �Uwd}J��F ��+�y��l{�5~3ڃ|�@�����}DŸ�37��xg�P�Z���)C ��F�l��hƊ�pԤŷ����+G���3��)Vy0�e>������s?��[��\�HL���T��Y�m�pM�ā������v�?/��C��%��Z3���[��I���s���m�E����ɦ��	����X�c_���\P��®�W�-,���(8��u�ȶ���Uu.��4Wv�8I� MY0�#�=�K�_BH:��%���y�d�8��)���R��6��������t�'�@������æ�b��Rf��̦dTr�J�.�8�8{�IeI���e�����l��ʿU�~��d{���DiwJ���杹�1*�h���������cep|�� c�W�̖�����xd?&�9*�{��C&�K��p�PȚ�M����wQ�eK��T��"�(
��dq�����R�V�����;��|~����+���`0���J�m��(=O���6ac����E�B+:��桠'�����O����jw_W����r���SZ���dcm�:�Ҭ�4�-p�G�GMҼ�Bjwf�7�y��2�����#��L�t[�`'w��}�3n�v�!����'���MM�aqH�xO�`�YC�DUī�.p5�k�K�Z�&���A^��SJ9��m�6#v�W��Ƿ�ÃU+�@����]g����E�n����f�����C|��!���Et�d�e�ŧ�gIB����=�E���H��L�����,��њON���Uͭ�,�]�4�	��9�g���*\�3L�x�H/7���0@pW��hƘN@�����Ɵ����/����?lPa��?����¾j{u��=~�2�
��}n��n��u�Э^?���,pQ���{S�D�Ϊ�˜�$߫ܮ)�ە�bF=��I��>X6>b��uK��ʉK-hr�� ^QKcN֎��3��5�}T��XY��K�6gE^����S��ZRje���%8^d�1�B"r��R;�v�q�M�!��k�<�q|�(݂7 �j��ؕ��%��*[����3�mk�B�Ԟ��T�g���!nD=�dI=}t�Fo"P��i������G8 �\ʂ�ӥf����!�۶E:�z$ ����l��6Ɔ���"��噣4{��=��#�����kt���T�-aP�j��5�*B��Y��
�ogb�aQu^)�x�C4ko_�
�}Ϛ�Y�)m��f���0���N�԰o:c=�s��@�q�v��d� ����n�w*��U֚��s����B9�cByXH}8_�R���<Z�k(�CAK�`���L��2�� ��>��)���N �x�Q
�vڳ��C����֬�3��~[�����']��~��E��y�&�b�O�SV�a�&Կ�]�9�Y5�#�� �3�p"�s �:r��,�	#� �����CՖӜ6�u	�b94���`�q�pjf�u�5��-����y7�O�|`��.���+�T��������g�rF4�Om��~��]�]o�Q�Qw��_��TH�������'��F�nu��l앆Œ��;�
F�t����H�kd@��A�ܵ����K(�/(7�牗E�� ���C���$����W���#0��{�sUm�t����C�M}��z����6�S��ސ�C����D�z}�f�EY��S's_ �c��"tu��$F�<��V�}e��;'��_��Dj��]��jIN�؁a�M�%�|m��@��}��M�3����%���k½%Z�gf�^�m�Z꠪�?�E����=7V�o�`	��I3|�\�0�C�֗TQ�$�\����+9��*`]r\��v$]��':h�G,��?U�'�P��O��k_�{u���YNn�07�����3װ��B'd����x��xz�iԢZ#�*�ݟJ��I�U��#Y��F�Ϣ�R!]�W��_�y��"p���REO��c�6�����)�1a2�@6G�j��Tт V��7V�QҶqꞋ{��wRI������Ng������B���ĸ�R ��8� +5VjQ�����<Iգ7����{����^�܏6� o�%$�<��W���X��
�]�8�KU�/֔9�;U�p��ﱀ�_;z=�������
\��ζ���P�aC�6T����i���'�?�N����A&S5�9*�Vo���ثs��/g����9ȭ lhi��mL���W�=����G�p�X����_��"�)�"��s4d��5^tn�%�������d�%�αC����x�6U�(`Wf�q8Ee�R9��x��z�d3J����S8�_c2 W�$�Ïb�5w��{�|���VXZ?��4-�I^�R*��%֮N�7�uj���O������ك�LR�e{��ߩ�H��Sl��'b�|���Ѿ���^�?�6�[��۝$`"��� �����vb���HT�_�@0��/����&p��^�[_�l���"��Y���klL-G��=iK�+�Y��+���/ �`�t:�G�.�V���\��L6[�-3�qH�s+k���e�T�󰶞B���UϞ�e�9ۗ\��H�z��� _QO����$:�{�}�����m��-~� ԾӦ��隋x�]z�:�Ia[�d3�=��T�����
��^*˶�����؅2��[���q�U�L�S�`��V�|�aZ�詡��?��>"t ͜ǛW��FF�\@~ڑ�4
@mi���&�:n��8<>�#�x���/£s4wQ��T�(��M��9�@U/F��ޱq7�Ϗ0�OXE��H�)�}�4��g�ۛ@�&(q�x|��7�
K��*�)�=,�or����"Uu�4�AK^�wjN����@\r�I�����G*��}��*qreU����p铙�8R�aE����y����h��#�5��4Hr��l��Ɪ!���W9~�OR�Ѩ7��Vy��9q����а�UH|�̚ڃ�Iɰ�&�"$�1XקI�wڿv��إٱt׺��(��P���hMĕ'�p/ǘ��s�p%�am���b�
}��β�j�#aDuJ)��>��[
:�ѝ ����-��u0 �趝y�\�o,���QVl�OXf�E�h��x�l�?븆�/-��p"b�'gL����b�S�O2��m������lY�i�B� �a.�>�
��9.�7�]��Zࢮ4���NؼV����k3�v�ny�u��M�}1�Tǟ���}���������ȿ~0lLM�!�?���y��M�?N>@��A��������@,�?� ߾��Y�V��n�> �)���|�I�|��k���7� ��[���"�~{����o �<�^�!S��`N�6j窔>�s�os�B�#��y��G����KP6O2eo~DxJ����U�p.��T�������@�&>�Q�9��Yg�"��>��ǢHuJ�J̋5��p�7A�4�-NE�tߒiq#��?�i��_ᤩ>��҇�������b��'+M4"��c���c������n9/V���a�sHj�wF*�bė 
�����z#��z'7����ա�G�E��Pe��`U����X���7'S1��G������n~U[��[�/��|���)]�fv*3;0��M<Dؒ����5kM����8%{Ō��Q������cC
��}�O	L\-���cL��©��:������y�"����;t�23X[�J���o���	��Vx�IV����;䟒V苨�eM�{K���pa��A
a��ª]|Q4������	��T^7쩤�5��6�4�=��n�I&�	�^��"CE���)�K�[H	.�~,X3tϢ�h�B�)�q�ѕ=
��.�e �o	<�2�rD2�l���_cQy`^5}�1y,'�� �q� �N�����R���B�@��iEH��VG_�����""�d�s�)�ͼ����1�+U g�ȤOk��9 ��M��<����J�����{�qPNpѩ�Vmx�ĴVHj�^U���Z%�G��Z�n0'�\4���^�������W��~����էV��7U����M�oTU9��: ��I�i�>*�6@��������ړ�4^��P�\�e<ON�Ka�� �B�>^z2�	�+�~r�^�]1�N����H*=��,���+��L��I-"�����|�n�|�Sv듘^���d��T��������_`��)��>�~�[�%]>ğ�,<�4��Tp7I�n8�l�X�<L�\���(���*EE��)	��T�^��X�?KLY<�#R������:�������Q�9A��I�4x�F���a�g ���-�P���p����Aj����'D���դ%&`#Tx���W��f�j��`���'�јC,��b|V,�
@]���!�������s��+�}�	��?&%����u����ZK`��V��Tg�������F$Rc|����Qz�^���<>W�=�֨��J�v�K"8� ��4/�|�H��ML��	Y.�^�/�F����J��>��׼�'����^��D�I��̗��Wn�*���n�J��#����~��YڀJ���b��^X�Pk.���%;2Vd���`1��ܳ�� ��
����<]P	�j��I��S�<5qΑd;>��.KC��Y�H�����ڌ����[ s�z�c���!鄬�[���8��WYe��o��	�=?3w�󣸲��<�R%}QMRN��B�"U��1Z�1\�-�*^��ݥ���A,�Roc&��ݭ���A�G^�'�>�4�jtn�dC��Il��ءg�nێ������U��C���
��9�pbQ�Z��6�H�]��e��E�w-J�)*��Y�|�<�����Y	�}V�JY�w$.�� Ty�|�ͻͶ<= )C#_#2����4�4q��[���,���XcU��x� ��5�.[��8�p�8+�j)v�.S����>�����-J.
���T�.±�6���0Bex���%�i�p��eh�u��j6G���C-�Mz%�օ���������_.%b~�(�'�(euDk�]1l��	�ǎ/JčYN��@U�5��䳳����C�E��t2�hB��}�z���n�`�9���5����ư�ԋd2P]����ì�qM�x�:Z|���ꪡ��4w�vB6�QAn[�*�"$!qɾ��I��< v�S��,Ծ-�j��xv}�!�:Q��$6�3�T'LΕ^򇛦������X7C���$|-�M$��֕�7˵4ۑv#�/��"������s�ٍ=
�[Z���>����X��
z������j�ꕳ���/<�ڥ�roG	��"��u��s���L�� c��p�sR0����Mq�KL�O�G���R��T�7�F/� \��SԄ��!`�|nK-�
a�"�4���k�9��!��/W䢊)��5��.J�c�����c�V͍���ƿ����D�?AમȐ�fj�F��F��+�#�'B33�~ʥI�yҳkt����5��let��\���9ޔ�bo�9m��ǽ����#q�ȼ�D0���M������B�1�9Q���p>��;� }��lR�w9Ӷ2TZ��58^#pN~���$�X��1��M�۠�w94�<{��@���^h1ןO�]��������!��^�U�۾�9P�`�V0,��2F��xoT
tOmq�>䮯��N1���չv�2��&	�?�m����?-lOے@#X�X:y�-A4��@���^(��xzs���2� �Wd������ci�l�F��������⫑�3��ӊ�cF#R��8�C1�=�X��R`0Eص�K%� 	��:�Q�)A)Gc�]�)Hd@+��WA#A�Y���"3�S��w�r�(��1�9,J�d�>,�����hz�����,�W�X��uU�p>�1���+M7�(�&�i�'I�Q���m�
� �9�0[P�
?�]����N�m�ɭ����M��ĉ�O��ro��C͊��0�`�ژ�p��N�<��^T�����Cw2����.��7�[��!�w)��&�no]x���i�f��l$W�䯎� K��(z������N�����^� \�j2�⺈t��RAfKU0�G�0L��kV���d#',(�	-5ځxZ�#���((>0��9D����b�rߓ�<�jsD|�构�6��fW!��;<�F@*m���v�O/'Q6E.�6���c��QC��>1��#=N��Qf$?��N�\�60�|l��k��,BC�rT��T7�C��!~	�i�żdr�//X��6�9>�c��q�e���*ா9�Y�C9?�I�A����:`7�G�7X�V������&+a��D�̀�E92��}������hP������9�;:_o:aõH������D����]�}�Wt��*)QvIK_��Fj�����gEG�����AI�s28�+H�`���:����L�ƀvm��ƾFtXl5�M�{[w�5.0f�,���tpާ�Y��-�Y��U��x�z0�r�u�U%�c{*C��t;S
�P78F����+�P�A{f��?�8 �&e��-�%f�_�8`�g|��H�'��j	]��O٨��Y
`�G�ߗ�#],S9��ͬ)���U�N�UR*$\1��T���Y�G�g�i)�����gfť�
`����h%n����cN����}zZ�hT�V����d��@�<�;�x���k:ț���w���S��}~e�d9�\�3&s��.��51�F1���w%��S3`/>��]=��Pҽ�7�������Hr@��v�U&P�>��T��O0�'C��#,`�wto6�K��["���g��,@�����1���z����%�QN	������'�����գ�>�� Lͼ��
�T%^�z/��&��ӏ���,u�~]0��.�]ZN$d��dFL&�(�䜞V:�`+�/��8��Kn���u���d�q�b&,�KZZ�K�۾4�r&��vZ�N�bT^��a}����' n`�Ӡ��.��b���m����oJ��21:b?iv�v�#8)K32�����"�hJ;	3���{]��-��%�Ε"�(e���Վ�>�\ֈ��W���x�-6G����2�Ai9n�UͤOp,�<�H7pc��W�K8���ٱ�����a*�\56��ል��'�?�H3���K:6s�g+(܅e{�Ѱ�V̌�������m`!�:W�3�����G� �̧-ub�u�o�>�gF�%���1|�WhB�hD9����C��(Y�p)��_5��Y�!㕌p�����=f\���!�g���zh};;��L�Ԩ��hwd������#(o�<�~k�ڣV,��6�fe=�0�Y�uTa�bq���۾َƿW(;i���fbױZ�^�D�Ԟҁ$�:{>�%�[�Q#�9
���>_�`n��!�yK�/C�H9�N��D���s+>w9�thr�t�J]8����Y����~��av���~PSk��fMo$� �r��q<���i�҆�@�ջ��O��D���@U����^=��Rk}���6�IC*��B�����Q�`6�SjFe��t�LXF��ӣ��S���7��d(�|���C0����}�N�O
��x��c��t�Y�6�����8N�es;J�8
��;��$���w�i$�	���Mq:O8�v��y?d$`Sׯ �{�K��TZ�)ur��ż�,P=D��K��Z��_Zҁ�&О�i�h�?#��􊘦{)��/�T�<W�ճW�.�"H���}�rQ.iX��sK�� ���,^�pz� ϯ�r}�Sq�d�\ä�{<}�~����1\��%rG�CAP}�Oa�{z�nf�ы?��I/rK�<Ŝ��E���& �ů$1�ڝ�Lf�k$]gH6�
�)������������^S�\��#(�#q���ƒ����N{y�lg+�����ڏVa��W��!.D���^�_�}��a�c ~-t�
� �,@-��9���k��z�ҝ�a�K�jA[2�QH�kk;�޺�b�,ߓ�(����ӓ �o�.�~z�B\�!b⭷N׊�y�T���CO�Mr�n����FЬ5r�~�}F�9��mL��J� ��j�f j��>�Q	]�l*B|�u'�k�~�1�:Һͩ��6�����6Y��h7�Bi�lD:��.���{=���Ֆ�5����¬\@��^��<�e	���t"f����}/���݉� `��eFl]L�@)M�mF�o����ˢ\k� 1�H 1���%�����w�{~8�ܯ���:��c��$r�U��48	�T�^�2~�L��y[����w�2���	�e�����dg�&�z�)��fI9��Щ��ia��o�G���m�� �ts��̙�
����-�D��_�S$�����캸&��<���\�:�*�f�z�"S��J&�~b�J�sڳP���7�&�~���L�!P�Q�{v�{!��6.Н�ڣ��c)c��Kc �2ͷ:����ur���![ʇF�*+{��©���_ü������#-�M+X�QB�[��m;#�f�����Ƽ:z2�;j��!4"	��:懫	��������Kl�B�i)2^��y�s� �6����,où&���
��g�K
Y�_��K��ޅ�ѹG��n��?��d�*\�(Ht
�s�<ع�^?�!2�Nj��(�&�>䳻��>�l�ܨ��Ґ�pٳ�#��x"�<r@��I6�qj�ߚa���At���"7��5���?x�TU#�M]��7f3����=3��JG�0v�ۆT~��5�O�gG����i�w�B(/��a�U��>y�OA��P�PU��q��j#���}����X��h�i��7�iR�����TF�)6���E���!����y�3�}b.���(�c�xug�k�ih(<�V����{I�a(~ �<��N�ŴQ$r��T��m{�&VM䐏K �
8NKdK�I�<����ŭ���,Qw	>���O�:m_	��o�����'���R���mu@����-ߝOL����gb�9/�O��J��o�c��/�D���k+zɾ���3�]�HiE~Ic#R^$eM�R�{��7?a8x�ԟ�[�W8ĜRJ>]��M$Clx^f, zI`,is>��ƹ4:���Ox��л63��'oDGR�"w�ݥ�&��2Cl5G���)�a��џ&}��_��جxf4��6Akl�ݳ)����p��#Ny�J����B>����1��@he,��N؎v�����	���8����6 F������_>�#R�n��)� �f��� �sW�9���ñ��nF��1s��Մ��x5;"Vzc'^��Є"z��כf��L���W����kia����_Q		���?T���*v�������G������a� \�8��=��P�'�	��ܻ^�tD��oNbr�}�4�yɇ�����8UP�8I�Lw�Hҙ"�.�_z�0!���Ɗ�j��ص���U���{^��-ژH��-*��K�ܦ���s��
/}�3X�4x[a�E$�G�X�}�~q�L�71�������� �Zn¡X9��p�]]���}��J ��]�}:�î炗&���>�QmӘ���L��Ι�������v��YW����
��y��
�w�����#�-��$v��k��e���m�8uw�f����cN��|d��du��5\����jR�!%*�i���KI�Gi۝��޳����z5�0����Vg��N�6���n�`=�	q�z�@n�(7`r���$�:���1��J�U�bc�a���3!�)�j�wA��� 7������i��_������1Ɵ��.�(�O�F�a1(��l�����l��R}�&*q�[&��~*uL���T�IܒĎ���?����4k+X�~�0����NB��޼xX����'�z�MVD�n-���9@"@Sz� �o���-W�C$5/o��I�]^�l�'n2gLf We�4w=#�q�����;'j��^!�+
��S�,�i2�|���\~7�RQ/����匃����?�N��5,�{8ѡ h�M��%A ]�8M+��"�ӊ;+Ѵ�&����Xԛ}��i�e�`6�FN����-�#b��@:���Ƙ"�-{�clsM��߭CR�١�J�2�A�L��Sb����k��J4��E�e�42����G���$b"I҇�ȋ>1ʃ,Y��I����Lq��gS󓏠/_���.�Ȇ�����>��?K���[Ņ#���/K��U�U�)�tW�����OE�L���3��ި��5s,(�2~�F-�]�[,�u�9͝���r�Ã+n�<4q#��t�t�Y�k�E"m�I�=rG��q,l�l�>��yp�-�^�)q1/?a��d��0sK���%88�RI�5o�����t�!ՊLe����)�ZV�L�aN�Ī�����5(=ߛ��7��!��p�~'L��r��2.��[[��J�rN�6EOU\�tD�K���}&�C�H����u)�?�M����e��/ �Ʋ\q�Y,v���q��D��)J��j-�C>(�@��5ێ�	�pX�Y��J��Ϻ���Z������gk�tyg�.2=}���p=>���9b�x�Bt�0��<y��%N�scu�������-���!5�lK��q�&?0�#̭oɖ;%	ސ�U�~�:U��Fj��y�}�ƪ{»o�~��<A�G|�u�/�%	i�ƀ0�b�t�w��0�3������E� ���L���}�Y
x�?=���\w�0O73� ����#Ń?dM���8e������!��ka���yؒ�wS7�e�q�*"٦U9�_�naQ��$��Z �TJ�iR����Ɠ�n�*��I��+v ���M�tp�7T1㜜�jrKjz-�akp_9���( q@D�B4_-�Z���IKD=�9�R�ŃDs��!D&���M̍d���⬥�Lϵf?:U�95ͣ*�Y��_<ƽa���Ԗ���J����|�$�E��>R�Y�	{jt!
���6���1���Oa|����c�dsl�ap�D'����!!�0��|���2C�C^E"����9�aP�gY��܉Q�jB[afܠ�(������H��2(șE)�������9 }j��S� ��{���@lTE9��Ǌ��g�8�9�O���A,�앥�-���t`/��w��N�uRf��zV�|��Y+�6�I�Nn�v��>��/f��y�:�#bp������ݦ=j�G��1-J�����1q�2
Q�[�b�­W��m�R�t;&&�Ӝ�����&�z�SVy8�d��6�
����BU^1�e�n�D.������-�:�v�x�Jʡ{ ��`�1<}24q.u)��w4�W�'�B���ݷ��@/p�AV��Ag�?�.�1��z⊐' ����ax���	�4$ÅϺ����(~y��:b�%g�fg��Nh}Z&w��Yna�*W�������T���
��AU����Eč��=SY|��p/x3�J������<1���&c�/ˉ 3�쪟j��*��^ʃ�$�-,1�D��&:w��#%��
�Q��\�m���/g����'�3�����#;�bS�6A�x��I�K�>�G�h���wF+A4G�خ��c�b�*�7����"�I���6��!eS��M����k��-�>E��+�{>�̤��:9ů ��������*��vpqQ�#Ֆ�����p܍ZE�S��1�������܋��@�F�3q�4hK�$,>)��M�D���a���=>Z�rܑr�i{Z�� ���������:�r;�G�`~���WAP��%�q�C�g��E�n�{h�Z�������U�Ym�@[>�5?8�hU�&��]��rF�_QY����p��d��3�k7 ?d��3r�3Kmq��Y��W�˵s�`]"���:����)�'�L��g;⯂a�B1>$V�9�d�v1�� _K�����+�29ңk��-�(�)�s��%�mމ����"\Q�8(�M'*�K�f���d8nm_�gyg/.7��|�E�q�Q�3l�����]����婃�u�nWn��P�]0���W�k`�p�<'�H�b-�B�����ke_��&�x���ɣ���>��M}"{)I�}y�F��3�z� a��Q��y�?�Zs'$ ����2Z�tՑ���=ۣ։>��}���*^�7���W�Q�#x]3wf���Q�����|"a"5����
"��rU-Ύ���s�8��J��E��t�UJ���$���S'����5���@�3��xs����k���r+<�U��2\J��>4�@�-�|�ʡ�o����[�ҵ�n���UI(���Z� ���X$�oH$YGna-_�.���2l`���{���&���ȋ^) s�$���m���_1fZz]���Z>��GUz�f*���7���Ȩ���M��l4\��0���@���R��"(4���â�[:(�>o1י#bs��]b�k�7A�)�C23�M�W,O�
�|!H�e��~!)tOP:$v2�/�S�=�O�f������iip��d%+;��:
B�j8k'�\�i�hzҸ����_��#E+�c'&Gޡ�q]�;[�;�iS>�,$�vs\��}�@g+��Q�rr�FO
ez�y�P�f.8w���K}	�N~?�?�HeXyg+$	SK��*���/��Ly�.���ml�2�'ST����9��A�{jJ2�%n�$��hb��ی��	��A�Y��i�����AG�{�)tg��Աi���d'>-(�2�\�J�\�2g�Թ�,��`ޘ�`v�3��Z��r(b�ƮeJí']MgI���}C���q��j����R\�6�,!`��Е..L��˖z�`��=
��G�Ǳ���������'Į	�R�6ï�fS��?у�:^��ʇc!�1��'������x���M�K6R����rI�>v.ߐt/
٢�����}7ϝok��y��h�,m8!kD/s]Q_>�[v.�l�p	4��q�� \5��٠����V�?ڴe.�Sq�[;_�O鏈R��c�CS^��f8��C>V_��gטv� �:gc"�G'���k��%i_���`��
Q1�)�V�T055�04�I�s`)E�@7d�W{�z����E�/�=�"��7��Ya�{���@W�SS�~��i�p1\�}�Z)�a�0�W��y����<(ջ%�s���� ���ß�-�m��5tK����fo����p��=���4K*Tw3�/y�_z�ka!�{L�X�E��ds�VV� ��Y{/of
�$e}V�����=W��9U䙊�	Ȼ�-xKðK �;kؕW^���v�Ж�|��,��k�ّ��-/D<�eL�6���*\\מ@���9|YB�P�L]����l-ȓ����=b��:�je�jD��+RD����W��95�����P�r�A}߀ڍ��d�ϳ|ѹ�e�	����񄌪Wؾ,C�����oY�m�6L�3�a�gF�S:�ʳ�x"p\�=�ЗOk1 ��] �%�{o�=(��ޔbX��E�=���{0H�������,�� ��T�*��"q�t.}�!}qB��	ʆ6�����{o	C�~/*4l����v�K>cʤv�RNG�c������t�g��gO���{M�Х0���J�y�����N�~�Ct��D��}�� �	�S�r$�T'�}]kˤ/�����2\��C��e%f�ICE�=�,x�_3�����$n@�6��\���)�_y�_~a���ˉ��ႎ/-���x�Y�M�!�]�[>�|l�L� �T�����D��{%���(�*����9��  �2n�i�L��2�-u����
��*k6���d�y/�nv�[T�|4A,��8V��@q�i��c�M�Κ����P	�B&-��BoWB�'!K���h�:�<�̎�*w����A?R�<h��F���b�B�}�n� ���p w��ON"S�e~���Q;�#�ӻȷZ~nė��a��k�O������S�r~�	?��&m��5c�	��Vz≿�@ICv��l*���Sr�\P=���NԾu��R�Ǎ�U���ԙ�&^��Ms�?fn�.�3����^���Y��2yl�$��	���˸	�GL.(<)��4��W��~����.�����8 ������*�L�F�N&N���� 5�X������ ��&	w��+�<�����O(�9��g ���e�u����y�κ�\Xٗ����)�Bh��ym����_��b*��_6vѸ�Zx�����D{�/���"T���Pϝv�,��q>k�qp,��\�q&.�����ܬӗ��>�/�1E-����lÑ�|+���2{�O�`�r���vw�k��6���P6������h��>e������}�<<F����{:!�ծs��@����s��^C��w\W�2n���j�oY w�w��Z��Z�ü�3Ͳj���a�v�Ix17�&�(��M#�k����+]���k�n�ᾌMFi뷪Ld�yidǦ�� o�J�.]��Ⱥk��xJ��.��<_��\�Zn��������[��HH�_��E.�PM>�&W��ER����mB��P�5�Η�.3��ߋm�gK P�o�?��`��1���\8ՇG�����j��2n�Vf���5a2"H�zN�Ծ����@P����1,�I�_G�`��jF�L��w�fa�5����ro�a챔�����~�4��]|h%$�U�$mfR,x�F��6�X��G���K5�*[^�g���9~}snp�e.J2�쁆�x�����coX��Rd��]��|�'}��m5�d�Ó휛��jK���
��L���<�M�֣2DĴ=����!�,xD�_u�"o�-G�C�CD���ez�JB���W�_�����)]̍^�	yр!W#:J��9IN���d�b$�58�Jm�w1ɘ	�~	}&�ݾ��� �b���g�����N�CM�����CS��0��z�gv���ְ��%P�4���kʳx�ik��%}�	��6.����>~�hw�/����+X'0�:����:V�H���h1D�8%���I1y��\7~����Ѱ�?j�VlN�^�W�]jB�4T|�`�P+�T1�3`f$��ŗ��U���00��&���+ϑ��f!ӹ����x�!���L}�ss� :������;(��"o�G�s�r[X���
t�b��;m:V���"w.��Tbѳ��*R|<ok��*�TU4��AW0�?Y��3�9Q����!��:+?��b~�ʮ-'f"�����;�soB�9�Ƕß9�Q�(Aɥb�ݲ���/��o
1�Ý��gPyS��T��[�f"G��>-�1g��5��6"����C�;����'!�H��0�vǎ�V�D�*�� ���N�jS���5�5r�J���8��Ԅ�V#?Һ��a �]���i}�������T�h��?6D� �e���*�]n�ެ���D��zW�:��]�8*(���̇���u;�.��
���W:=��Di)�
�I��\�s"W4� i�[��3����!�� ��o���<�_]��6�����`�nu�=5���;�A�f'������0�[Ҡ4P�� �9�E��KO[AO�n�a��A|������EKS�Q�)R�	����������M�7r����l#��%0��|��{7�t�Ѩ�V�B��d�PYB`���k|]�^�(S@�K�N�)�\�*���#�'��d�����]�0Cq���gN�����J&gu�0q����e�b����2�Ǹ����s+�s#A7LB���2��j���q�˚r���X��M�����3)��]�!Rמu���
�͏� f2�蕔��O��a2\��^p�b�����L�,y1Ty�L� q��-(�v��Ic@K���5G$W�Ԅʜ�>5b_�����h������@yCt_>�hÐ*�r�kS�
��p���4Y��c��'}e\g���`�ϝ=!� 1�4)ɯO�Jo�6qN�~�`��Li0P�������ݬ���C����kD	D�&��sm9B҂���xD�)8��y���ڇ��<��v�x��W$'쪙�v{4#r�E���=�x�]1��5�u"JD�6����U�C����T�c|�(! r��q4Y�Y.�S/�)Y��Љ�? -�v�	0Og�T���ɢ�r8���qfWUH�J�z��_҂甭�(R�9_0��M쭌iA��bY�/fnr�C���uϹ��_�S��A������w������H��+e'!��
���`��5BZ���ݬX�����PP(ۆ�x��^֩C�h,a"�v�Z��5!�.�}S�*gT�^͗����6|�v�Q=sY��֧�c���"i���*ϭ�P~�(����J���z���Hj�pi�Yt�<g(C����C3��]������F�!"*���2�9��a�Ƿ�[�&��D���D�e=�y�5
s[Q�1�n{Uڧ�c?�ߧ57n�P�oe.��#���Tb��0���N�~��_�<���s̛��ɋqY6N����[��st�ڰL��t�R��wl��F?A��No�;+�Y��lL��#B��UH"��dB2z��kdt���H�Y>�4wd;�����^�gs�\ ���{m�v��l ���~C���M�S/tѰٱ��dUOR�Oԓ��EΞ��$���
�-��'w�&<��91[L�����WJۺ����R�� �� ����l��
q�:�;Oow�C't�~�I��n�[��R�yh����V�z�K�z�KW���f$G3͖��B�bOv/+!t��5����7{t9�7��G���!?=>@�^]7I�����F6��.�X�[�/{�Yv(=�Y��E���$����c8�ÀLi�O�v��F:X�G`�o����;Y� J���@�oR? �q�o�]=:��_����-A!t������l^��IϢ��+���k�����!����L,p|@gs�3D�9ׯ�ȟڿ8`kP�mm��|"� n�j�����V��F� �7J�PN�P�چ���a���VW(�����XP?%H]-6$+OZe��-Kq|8���KMk�-�11ޚ�"ƈ����~�G]sB�ÿ�D~��,3~P:F��S	�u��Y���/%-���� �sЫUX��u}u���]�m�U�i!��Zn�[#��0F����x�]f��8;W3N��cɕ�?�RcdᆁU@I+0�m�7٣-�z>q�HxH�ʋ�.�Y�m�'s�lM�bN������&�|����^0 ���+E�|������6:�����,äl7���J� ȯ ^ЧK~��Ƈ{*&S�R :��$�B�wq?"�����!��1�S)�5ױ��?�&i ݣ@���]g��lNL�8N�z�?ǜ�.�" v/5e`�i�3wT췍���H;w{t	�[��6�9�z2;�ȳp��8P`rX��Wh4`��EEĒ��1� �Af��/��� .�4��	m�d��C��Z�u,X�K#��BʝǛ䨪�bY�P_�.t�Ʒ5X�9��b]�ދ���&�H��謹00^u/���ʍ.3�O-�����~+�'^ʣv�d�MqJ�A�^f����pֵ��8ɇ�f~s�`��owOP��W�p8���� o/�:;����]@�<ߖA@�k��mș[�?�ӡ�b��{?��q���V�P������؜�4�>m��T$0gbd��@.��L��?���/#���[}�A����h6�S��S���)���Q!�g���^(���5��faug�����T5��`jP�^и�Ev��ƕ�;n���e�?8����*�)���
H��
t�Ѧ��=����9��#��ޞ|Wpo�&��_ 뗖z^҄�e7lQ#u�\>��ӈn"s��O�����w��2��W���:�1;�u���^�p�(��>9#������{��b�x�����%/�}���8K�s^4?q�"�v� '�J�
��>FbAj����/���bbqRuid?�Jk������9e��_J���n�5%[� ���ST3�����_��w��@�+�0�t�G�:�Qk�H_��P�g���8�8�ڑ�>s~���	��͆B�#V��]J����䯇j������;����K�B��=6�i��CRL�]���[����YQ��þ�UU���Y�y�U���K�������Ck�3b t�"	���_D<�-�� x�������Z߁&ݞ���KH����R8��gl�t.�*WcgU��۟��Q���ո�6=��N���׉hwR�❗1a���q��q�G�@��%�����k2�b����C�oY���Tj��E��h"`��ֿ����F�ZFa-X��
�¤��J��^B3��G�E7�ѵ�Yjf-宏�?���)^@�e�'�@CX�"�8�O��:BCm	Nmn'�n �IJ�W�C3a�_��ҢIF߃�+��ܜ˝0 F�%RD����Z�S���B�H"``蜔}85
O��f��Kd�,����v�0��\	4���d�ݖ�.m�_ ]�Kb�r����D{��s2>*f�:���)��椾(�A�mt�?0�`���(�^�%d_. ������Ĩ�ӑ���£�d@H���� v�@ �|��� �K��j�t��қ�d��{��m�y=-�Xg�A�l�%t����l,+"�#5��%K��jg�t�G�F r��p=�1$�3��A�r��e��_�Ƿe��nc8����(�DX.>=�$d���x����&�	݋*]�r̞�V���d���)R+F��;N��%��Đ�������d]��ti}d��:�QF�ŧ:[O��]�h�6��lX��fD-�9������>��uC���#(�����Sv���� |�F�O��)Sd�	r>� �G��j�|�M/ã\8�˟�QY��P�&iBsK�3�)���K	u9���ڞs�N�.Ή'2��"��v4)�������A��Z����!����n
�4�Ce�Md��F=�ׁl2ˠ�����jL��.i_���`��D�ff�g ��mf�8�Ԙ�x7�`U�`�諍���ztʏ7Ia��>^�_g̐���EAk��}��lr�"�ԙn��4gF�ب�H%��Y�������Q�DjMysk�їs��u�`���9	���_�����JW�;S���Ǎ�� np�c���:ԊJ�ƀ�Ոp�^�[!�ń���V�햒MT ��Av���[��cF?�)[>����&9݊E��%���¾I��֔;��Uy����b� JY��@ ������u/����ȴ�u�C���cPb}6u� J:)��k�I�d� ���D�F�]z)+�j9�W��� ����-������m�)⧷���e�c�S�&�r���\X�d�?��W�9<�k��!	b�Ӹ��U��b�ŉspU"���ت�mó�6�J{C�����9�R�^�������Z��3��t�B�Fij�8��1 Yl)���5'�.	_J��b�<�jZ���c98��pt�E�*�e��UG1q�?$S���2n������@�����=P�7��&򘐂�i%��w"�X��Y�q����Ri-����1"�ɋ�|��Г�����@�;0�IF�DX�h��90��[aO��!SQ�q2�hyPm�?�Yn� 1��ש���g���MF�'\y ������Zb����I���??p3a��4A�ؾ�m}�n /��CK硚��bj��C�uqW����tE���eg.�ʌ�#���JyǤ���0�oLb�D���S��}]���^3(iM�n��t�G���SW^ҶaI�J�ŭ0�H�����bp�T��p`���D�U�޴��?�q|�@'dl�W���?��b~�����o�̇�s>=r�3�؅��q�E��H��z��e~���7g�)�`�D�+�]�lx7Vq�����>�ʥ!��2�&|ܢ�<)�D*���g�͈ޙC
ʘo�P���ֶZs7"*B/��=����Y�/�>DGhӭaN� �,MXGR`���x��ÖL�]�}���A�6�* ���d�۝Z�� �Ki~�B�M-����a��{ ��e��e��;�3��Pw�C�*B=��N>�Z�t׾y�z���J����Mm6��v���ZY,z�0��_�m%/�.�Aи�]�ĥ��K7I�cU��'��n��J�(��R!����P�����2Iqm�p�Z騰��4�r(��{#P���'��uro���ju���1�&A�T]�� �"pb}"�F��Lq1ibƁ�(�{"U^c��ʒ��`Py;�y�ۣr؍���4P].{�AwԖ������8�π�;��.�n'v����:zd�56A��aI��ɭ�B0���m��HFw��H{Q�1�]��h���\z{�LPf��:��VY�r"&՚2�C�˺v\�Z�D�8Bdl_�:��S� �G�h����ե��/fؒ�����Ƽ��Uٚ�S�nd�tG=[�2�K�W��:@�(*���ŔP�=�Q���\�~C��/�������J�����IӀJ(�0�&���dc��"�vZFc�ƍ��,�2];�M������N���Z! ��	;��"�;b"t�6�Ky,�h݇�p���c�d-~�2���z���O���U��*7U��+��o�V��2�w�iS���t���*�[�����~�%��l
�
?>%TL�c�"��" G8V�>4π��N&0�f2/���*yB�L̺j9���1WWj����j�O]����u�zġ���9�$z���[am[�_&zP �E;hwL�z��o�����/\�2����.��ujQ�AO)y+a���nKR��ՠ�k},j�dra��[�j��8)���y@�`/����_tdF�3��Gz���M�_0tR�κO㖕���(O

�Ü��-G/��V����N?6��Ƈ�4�[�~!�C��9�+�c����Ľ&E�/��Ԃ�>��g#k�=�r9k�H�{���A���v8+���b.����q��	����=-�:�69�%)o�$ȓ ����e�(��#�=ʸ���Ɖ�IOj9WdЮ:xmq��4"�<�O�|�O�D�c���F�',���-=�D�n:�R^t�p�K�p��?�*�o'���H�����rB��6?�F�bs�$X�o����Ua���,��Au��>���R���S�4�j��>ü��/�������]U߳���ձ]6�׽�b_]�qK�Ľy���*�f����$��s�s����PS'��S�����Z���rⳕbAfm�%��J����cc�
���E���;�����������d>M��n����J���6ve�5�e����
X�]z%��r��p�!���K����'��?N(a���b��;��
��;k������`��h���n����$R<����|�a�Y��
��	�0�����0����v����́���t����3B��I~�1A�y��k��݄�$Z>��[q����!���Q�{r �K˟�Q�ϑ����5����AQ)�dğ+����d�������jr[%���3ݥpa$R�g'��r^;#�d4�=ދ��c��Y�5��Dbq�����u��l�A_����� �#9��xwH�ZrL͏�+
i&8���V�����<�t�e1�	�g��1����x���S��љ��Ϻ�z�#���XW�+�~~Y�j(�����j����c�����a�ɨ�ү�H��f��H��#��`Uk��n�)`��}*�0�ӽ���P��]��.�4�j����B�̢�l��ݏ�\c�ٻ��t���p��cO	\��G
A#���u_%�ҘD��jO5jULH:��ޯ��Z�'e�=�C
�uW���!j_�H��@م�6dʖ��l��#z�p��������Y�xӅ���,�W������_9�&s���ӏ����^�B��VV���mQ�@�{�t)(�7�=8m	ݺ���UĎ2
�ja�8���2x������.�=�e����&������ͥ�Y�9�ľ�,�[Wr�������,��o��Cj�vm��O3g)�i��>�/�@��q���Vd̽���C���%���PP��?�e4J
��}�9�J����+��.��������Va��������r�����&�XZQ�Y�!
-�*U���=G�_���HVzC��������v_�����U���K�����ѶlAM;a���}Rw�M�p4����+���&��)����W�\W��#5��˷S�QQ$Y ��R"��(f#huYCդt��7��D` ������$�m��� kɴ��y|������Ơ�K�����d��ד�Y���C�8ɴX�m6��%3P˺��Q[�tt
SwL<�ԩ���������N��]���C�i�̷�?��������?�"K�䔏v$k�,�� �0C/�~����m��lx����P�Hj�b��E*�+^��#5^Q��;4(z �v������ۃe�n�L�r@�-�pi��Y3J�rձ�wN1ٲ�fR51QǏ����x��9Y�)#>v��2�QWP�s���!z��E��N�K�㔜Z�����گ��US$l�G+I���ʃJ��[ȴ�}�O��E��W
����	���,aو���sF�&׎-f_����^�*� @������yI�ɫ�ADa����p��BAN;0��q��Γ��/�6��A�-D��%Z���Q�t������Bڧ��w���!�y�lM�@G�p)G��B�c�x�΃��GZ��U�����2Ć�����}b|<���l�?C��0dF0	�����S!�49׊ӁP�yWA���ˀ���ai�Ș$ۢ���ϭ�2:��%��'����K���2��*5��������8K>�����G���|c796*V��F 
��>�hJ����ӓf�5]宾�S�&��J�3K<$s[��҇�\�F8UC|�Ν(��K�C�#u'��8�e�5&
[�p 1U�����:;]Z�%�̔lk��{�jV$��G+43wGA�6��^}&���/�R��R��	��C�3��;���ӡ���d���c@;-�6+G��5��Q ��ױj�9H�b^I�|_���{��"�4=!��uUђ�0�WH��Ś�౫�[�n|�@��w����R�{,J��(���}���xѵ��l���7]�J~�M�~��eL����uM��jN�5�Kj6ͻ�׷�`c�%�rF�W� �`��k���Y�R�TW�w�o���{c�e0�֙zr�`��,{{O�Gpf \�u|K���d��;#��1��%M�H�Є����68�Cʅ�����2ԟvu���\b�]-Q�_j�{nr9�mUS}�N�h���hKO�hQ�e�S%'I�3�B���}��(���O�c��Εx�&ůO��];�ϠT6m*v�R�Y]�>dW�k!J���'�tO�)w�k-��}qג[QFc�~���%�����X���8!�V�?��~�������_���*���sPw�9��{�w��ѓ�{3ӣE���j����_�����/�9�*!K�����L"Ze�S��M��{0j����l#'Q���y�����m����1?����Q�PΏ�Z���=���S^#�~�Մ�y�w������*�R�F�坎0�۝%&��/��L���6{��m�{��G���'�v"���y&'n�p�;p�x�qե��ߍ2�޻���	�TqӒ�m����O��^W�Q��(�Fz~�b?�*~Ƞ��iΒ �JT�.eR_I�IY'L�%	���~��� v�J�g<�am��T�x��J����=m�?����%�͜z����C��aA.ф��Fe�k�E_�p���,3�Y�&%S�T�����i�7�R),���P�7t���M5�����x�d;�YU(���*j��t'+��C�x���Y�pn���.�>��'#X�1Q�A�� D��0i(Y��%�`a�쬟G��U���塛'�!�\�"R����s߹=P�%��g�^�m�F�󆨷R�&�x
a��M�(ݷ���%��*��s���L}:1K�x��w$b�j�T$h���Ks�8�A�P��U��E�W���ljS�p�%�|��Ţ'PD�c��(�b��|���`;ӆ���(�<�Z��,���7X,-��obQ<)����9iy�q�+:���^���ϡ(L#Q�Ȧ�L��O
�m蹐����KSy�0F����z�ֆ(=�d�ox ����F�� ��Ȟ���6�iQ0���F�e��l�>�l��K��҃9��J���a�����։��c	�Ďb2,�u��!;�ɶux�a��)oŰW�@��pL��4��?c��%e�B�\�>.1��1ߣK�\Ƽ|���e�zh!�-��B��QBǠ�7!��@h�>��7}y�'�95�����3�ϸ���L�c�#�!Ν�	����k�W�Q"A�"+6h����'���u����ӡ�<�����2J�ө��6��F�g��Y'���b����ng�ǝAXӀ��Jw�2���z��h��6��ݱ�L�r��v�u��{�_���U���h�K�-���,����F�4'�%}��c�)-���g-j��Rz��z�?� 4	ʹ_ig9)�����J>Y �?��c�bV[qb����J �(��!�J�ە]A[ǭ����|���Dk��	�������5gɶL��Hq-Ʉ��tv/�5��.�M����^���y��J*~��߇r����~�DA��w��?��[�!��K�a�wMuP�[x�"�v��=�@�Q���]���]�`���fP�a'�4M2���O���@�	�' �I�a�\3�5�O�'4�2������j�֘����s�pZ��$'�Ϻ�����?�0w�O�tT����m0cY�XZN����^�H'�z[���?U1ۛ��d��6�\�}���HdB4-��qb�#K������(a������cj��6��9���#�:[2^�����xI�"�Ջ�s"��m&(��n�b��ݗ�$i�u,u���U,~�b˚�3�^����j`�{��'�D�9o�\CoE�_�����l�y��#3as	�Q���"�1:���r�����~zi���YV�T3e/U�j��.���Ыz_֊@e%�cs�B�Ф�(�v��4yM,6V��F}(m�Q���&D�xM�0��Th��okʔ7&@���\́��p9GQ�8�C��`_ X���,Дq�Ѩ�2k��g\q'�rE) 9��	ev?�ѻ��P��g�"��X&�����mL@����q
�����b?���gz�b{��l�bZ��+1�����'2�%p]�5�G��:@�]���y6x/�+��б�������s�){懧�#�~��:X'b;���������]P����_��^�I2��{�U	�CnAeuyt�y�[N�Mz4UfN�3�ڍl<���틱6	9���ן߃]���m�������C�)�򞯰yP>�^Z9��A�sx^����H5���!���w� U_>?�(L�{Ov���'b{;����Q�x��dm\5��W���5�Ƒ�5�A?�c��*��~�����U"�Eq���eD�Z�}���b+f�c>eб��Lk�iSL��(��b�s�bț�d���ueEg2�;>��(7w�:����ڪ���k�狄�08��i�	)L�؏�w�
����;�G��첫��q���H���|cm%�/��T��r�޶�>]m�a�����������1�z>��J8<�J~u�Cs2y�п�����Bi���/Ĵ����2�B:_�I��s�k~S;�v�0�c�&Z�t πє��U��6Q� ��nn�����0b�Z'_Z�8��#�綫㘓��9'�=s�����?���_��e	�ZR��z�T�m)�*]�]v(��ah�Q$P}	�
7��ӪK�L�`m.7|޻a��S�#���	�$����X�K����*�M$��J@?t�$Բ��Iv�uQ0��ݯ-Z�h�B[�^f�w��Oy�Xý} T�h�1ՙ��\N6�/$T5,ߞQ%����ϝ6+�9a��{m1*@��Q�L]Q��q�x�[`��R��dȢ��,e���I@���d� ?$6��z��O��+:=��w<�Q�����mv�(Å/���ջ�}(�� 6��m7�5?���L�5���fj��8�k�hvhϘ���;ĭ/��\#G5q�;�ƍ�4k��^��
���v�o`��=R�����<������>g#Qì�W���MD��N��!��}#P���
i�

G!�n#*�7��g�R"�}b1��v0_���X{�ߑ�?���E��Y��ڂF��I�CtW��p4*OG��Cqy��
�
"�j>KJ�fmmB�FVn��zj#��#��Ĩ��iեl���_�Vy�D=�@��c���ڧ����y^��E6���:T�H�/���ñA�+����� Li�`��@q!�{x2/�=�� ����؃&�t�j
C���f0�HyZ�.(���rZ�����c�f���5�F��`ƿ���(ydAy`{�Ea ��W��BZN���w�� �Ǎ�=��g��g��	=`^F"���g�X��Gg�����7�-��=p8�5YXm�2�1	?����z;�������6��V�b�tȾ;�Φ��� 5,�]EEW@����[��	��[���[�"��O׍c�~�F���)�-���:0ɢ��_zʰFȡ���?��DRNg+��㑮�E2�M��+&�*ծ�<Z���m����֞���4'����H�%�2��I� 6��2�f�ϙf:r�1ͧ�"�ni�6�S��������Y}~�{�P0z�'A`2�=4���þ,�-�����.�����c�Dp�T�-��[��ߪ�%��M��o�p��f>q�U�Bfs�LrKks��M5�xI��I�;m0m�
X���]��z\;���[o;ꦁ��hjwM �j�ɟR�F��Vt���Β�]g�É
����P���h ���1�P24L�E���xК����������ӚCd�۶�D��g�{�m����V`1K�Cw��[���GpފRoB%Ũ��W��&~�%���kQ�O�mPo���!@� s����Q��Uٝ&}�7�R���{XMN��a�{)��Ƴ�j�EQm3"��U�3|ղ(o�Y��$�� ��dcU�1'�mu��z3&\n��S%Y\��P���g���]�L�{2�e��6�pT@}!/�?Z��HXe]H���T�$<��w�}SUt�
cV���.T�&?�ʰ{�_ݠ�@��9v������[����h���ul�@���lu�	��8���'�(��X �_���z܏PE�I�*���s$�ǃ2�=���y�`S#��n�6�Hg���_FN��i�7�~�T̓���5.��vs���eN����erX8N��k�4�a�{c;�T�o
��t�&�Y_���N�.rkbz3�����iTx��ŗ��aĄ�=r`* ȗ�T�6�.8$��ٳ�.&s���oA�ܬ���>ݬ��!�bW>�E�����彋�ù|[6C���ە�c�73���}u�6�v\}��J]�C�d�4^|�d�:�p`C�D�D���x�Q�nߨ�Pg��v�z�n|ւ����������3z��Y�+J�[9鳾&M��Y�֛�P��q�;��\�p�.�ߺ�l~���H�=�5"�$&�E�%���̛$�l8~0T��&<�AH9�H��L�I�S���Y3T��J���0��z%k�pt̖៴g�.�==����D�ĭi���PS9�g�K#�����x�rA��
�/+���78N�~�l��.�]0ƃ��vI}B5&�ןC����}��DzM�A�-������/eo�K��g� �c����,� �wF���Pt�T1'�$�b�(���psHh<�����S�9��:V춞ܸ/�w�P/����P
��[ݸ�D��"{o�`D���UZ����;mR���B�<-���}:|�z ���S�KD�>N���$� �) )��!���/�0�?(�����%.ƩI) ��8���#�'X�.���/̫�Xa<���Bŧ��"	��:�:A��rי@#
�?rS�$;�x��n-�*ȓ�2��nZF�,:���q��>QG� �.���߽�"^Z��]�۪I)[G�yMʬ��L���6�ux�3lCg%4���^%��nTC��kmd1p�2N�����0�,��5�FS6���.�-|�S�N#c��_j��eA���gٮ���NVB�g��L���L��p�kHw[�e�m���0)B9G,yD���'�D���wֻ�Y���ݥ�'��DmJ3MqJ�wq���/�k'� �rXZ��Q?3/z�y;�U�k�P��OԸ���ó�J�*�FX)�T@9Rnv����v�*I�`�"6�1z���J�d���/x�V�z�:<���]����F�%�>ꄌ)�xP��4J���w�ཌ&��v�@���</�q߯�z�YgL#)�׈�i�=6am������2�t�**��p{p��Q��김m�}	��(��FFLn�)�N6i�E")�d�*L#�I��̣�?m�}�Ж��c4~�Q��o"�{;RW��?��cZO�6kEJ�M���dg7=�֜*Ӊ�d^�C��(f�´ճ:1�B�xȍE͑���@����ۄ��m@jo��R!�';������P1�O��z�E�ٔ�,,k�3�견��������P��1���a�$�M��Xk��J/�|����:��������9��O��,���+��3�>���K��hࡨ��y��J��TZ.+���\�kp�����'���TC��LX��J�qMz)ː��Z-���&�j��Ξ�}�%e��6��o��7��������Ԯ}�Vi�P<`=3l?� �Mo��bo�!�;ػj����D��z�3[�z+}F
�^|�U*��r+Q��K~��q�;Z��'Bq7!���fʍ9(��w�t1�M��2���	�e%����R�&9��c�CT�� ���`�Vx�x�/ɗ����eHnEW��M�MM���'^&�� �Ŀ:;�U5Y�*�f06I�Z�T᱐^	���@aQ%���Q�ɺ~K����]`���)y���A��Ri
̧	)�W�J6b�?����˃+�5�1�\AIw��
}��~�Q��5����R�)�rk������Z�-����`(�����C��<,��Zo7h�@ˎ3j�|��xp����G�����j;�L�9٘~a���%��w�X�'.�u�1*�%�T��Y+�&@wA���7��|qh�Qu�Fcw;�m�2��7�l�)0ʪt4XԤ���XFW=u���A		P�!S��RfH�`��L���ryV��6�1�\����<*�yxp>�~��q������t�+;�K��[�F�������c(�z�a���)HB݆3�?�QF�Fv���a'�뾅�X('��:�[{�e�(`��i��?�`��o�H=.ҐizHu���\�K�Sk[��.�"D�I��	3���.Z�\p����q7�&��B���c��>AQM���pJ�<��Z*X�:�=�W���1�����kX���>�d�p���ǅK������],5�Mۊ<O�G���&x�h8l�#"=�-�$]Nͩ��Mؔr�y�B0kء8�O\D����\��������Ig�Y�VJο͘�.k;F���L^P�~�Qg��j��-�a�l��������5��o�3��5�����=b.��p����E�ә!u�������c��j�vG��.e��wg&RU����{B�Y�2j6�d_*�O��/lvYn} ���9�].b~���i?���&�浘I!���z��v�o[��e�zH�XSt��x4���]�p\��m�!��H����|�h*V��07회�S9p	Y�M��("��,_|<#m�h����P[I&�S��o�?����������}�!Ԋy�����'8Sx@�Ɩ����T���7� �6�7���^2+��Bd��FC[Ѻ(Zt����_��.��V:_��A#���4�u;� 6V����Ѥ���#������s��l}YO Ӿ����iI� �;��hoA���|��N��ְ���(r���o�7]m�i��.
�T�b��mE��~UõVIF���Y5#����ǔ���h�����H%�9Qjk�a�RS���_瀲�7�G�[��BrYC
�˭����7�I6��!
�c�?xq-�˭xQ�B�4����jM�wF�+⬒|��dѭ8��a��(Mرo�Eֻ���֬Riw?�w�2�E���2���Ϡu�7�gԜ���@=�(?B�Z�\O����~�b� D���y�W�Y�og�g"+
�Aރ��$1,ױDO���t���2��̇A����׾�w�Ů�� ��G��R~3��#I����9g�Bj��䭯 B��0%3q���ӫY
(s����R4%_�+�9���� ��%�x���u�α���WRm�pj'�=�ַK�b�_������(�
��W�-M谙�N肒@~���4?L��1nw3W���w��:��=�3aO�����������2z)��*i�5�w�.��~�	2�-�7���m�������P������4�kZd����u��L�����{8�é yS{���,+�i�f�i�>׵r��p��.��`�_O�L�y$ҟ��Ne@ΛE�:��	����u�:�����aL66�́	��Ӄ�K��s��@)l$���C�2'���ۊ�;��7�W���ȉ�<Q��<ef��kv4!X7�t�ˊ��E-X`M�����?6��C[��&L/�r�8B��WS2�^�5O�)�I���?h��rN�0��A�MG�\ǁ�@�,<u[K�����Ĳ�]���MCt��w�+�$gM$Mo���#Q
�ťv+�G��~T����]�Eh[� 8gԸ�ϙ^arh�DJ~��g�s�q�9y���r�>�,E�wJ���\��[��h��dv�i؍����UQ/8:o�&���H��%?���F�U�G�2�'E
�$�hrP�*V�zmUӯKؽ��܇�2���* �-�1V��x	̗��R3��wNL���@�
&[J�zH���;w�/��-�0Xs�Ӣ��ތ�t���_�)�|Y��'�a� 2@�F0'q1ж�P�U
��73�+.�&H��Ίy�[���b^d���������R���x�?dk���Xp�#�_?	j�'cC<��^F3u]Y�e�?�_<�n'F�`x¢Z���R(�M	�^��A�� @�.0�e�P[���`�L[�S=�A8
 ��Z�x��㜉���axs���ŜO�2Tr���U�;2S6Nx�NE�(�Q�� ���ݺ쫲���_��ho_��ҭ�7cY2N.�}
��b�/��3Y�ೕp#�-:x��f��YY�L��5�N�m�VKs�!n ���!��毧q�
�q��4.�#M��A�y�Ub�B/�Җ�ֆr]�{o���,5�����q$\;�әP�zy:�
��I)�|�\��c�%��=���'��		�^�Y�+F�V!8��ϱ�6�}v�m�`g򎙖��̒�i�� ܩ L�,a�i�����4�(���hn��0f/q<A�%'��n"�ڜ��+�i�����@H�}̻M�d_�ي���k�SL|����r@f:cQ{cX0]���9���΀�3�pk�� ��,����^�u�W(����������D���w۱��)���Z:��\<Ԃq3�q.���8;H�����T���L��"NM �E#μ<�(�#���I,Ч+~���k�â'0+݄\Ŕ�v`�mu��d`��Nm��Q����[�m��9'>�\�F�@��g��8��G����/��cZ�K�ƥ���8�r@pvIt�c1Kf:a1�o���^�Fb0y�Q�����(�
�G�2������`��k��x�,�w�\�s�y��k��ꛁ%��%��E���zd(K�#��X�SX���:#�mG�B�T�h���}M�˝�=	��L	\�ZF��_D��`6��cb��x���U��01� ��M����|{JK�X����3�D$T ��>Km��Tn����� d@�����+m���tb��0#"�3l���Ɣ�mLP؜U���w{dzs���61Ve��!��TL�r�3�l�v�Kc�.[�f�{c�w������%�];/1����*]LF�������90��]!Hq_E&��,R����{ZjI7�C+.RnF�/�j��lU���7<K"Q'0r�ln�'b�.S&�R0��=����>�U��$b���� ��ݠ���l�&��,ώF=�����R�}IX=�T)�%fX��{ŦT�D��~�����c3�7���y��tf�i#��7��
Z���eqv/5M�9��ڋ2����W4��ņZ"!ݤ+s"A��k�m!�X�=�I8Wp�k�ŵio����f[[;!�����Ģv��Պ=�j� ����bX�DR��0y��hȦ�����J��p��Εs)7����|O�����w�,55�s˒$��;K��q����G����騔N�"�v�哨u���?�m]['�&����1� ^�ሊ�-�URҘ�acf`�m!�$ظ?i�;�hm}8)�;��v}e�g7��Dg����=���婂�o�}��q�)o���Lzȱ�v?��&Yi��$��,�@+��QW��/$z7A	�s�|��BށE�5�
��HQL�[�VA)]=��ⵕl���uhS,Y���S���t �v���1���q�+��>]��ioT����ؒ�c���_"��TOW���Q;�K[�����UboP�զ�]�!lP1E_巸��57cOr;�$z2x�u�M;a3z/N	��"}������zGd��V����+ॆ1��D�\�ͤ���s��("�e�Ӂ�4Ç�91�R��Kˬ.�{G���q��A:���?��#�5�� K5��\LW�Ӿ�|(�::�J�fY�}��)�L�h�Ğ|�9��{�1�s��~� e�!μ���6�Cd��d�hρ�ق�n�(���7��>���~��Nv�':o���>��r}v�̓����>w2d���@RT��ۅ�vC�;F���,���JN��dz)F�.�^�؟�!���4]�C�"����͊iv.�C��oܩ�ʂ��p�
K��;�&vZ�N{��������Tb�`�����ě������6�P3ۼ}Z0ڑ���\u���?i4����(bL���y��:vG���^X�*}�M���6���'� �/{�K�dMP(����i�-�D� "#��e����Vq���X�7��Q�O)J�&a��W�}�O�x��Ρ!�ao��5K�q)�1��)��30�ʣ� �fF��,V�~�;N��>J0�}�	������}��-!������@,������b�}������g�n1�u���B)'�0���Yn@��%���^�Q�g�|d�o�}&����iJgV��/�;�3X|_�[4xMTU*��k�9T>��$����5���l��l>�2}�]G>����R�&ŏҒ�.��:|�1>������؝�1U6��^�f��H���̭ks!Cc#�E� �)���|dtݡo��Kz��X��2!���C���=g*�H]�M�~N�����S��4�ִA�橯GM�5�t ,�q`��2�I��2~�_�B��3-�Ni�	$��������
j��}�>���i�:���L*d�z�MT4{� {�Gn��ƒ�'8GX8nM��*���{�\���f���3(�aؒbX�wۄ���j�Fn�M!h��j�;`���:�ZH�of6@��' T�8׌�+١k��&�޽�8��O�+oke�}Q[]m�Y"*���G��a��`�e�(�D��L-��0UR���K�G�A�LM�Y=/4S3���T���r��R������4��U��%�Pid�S�%
Q܏a������~A/#x��	�)�暖�UԤ��D���&��6�������5�V�`�a�	��1�X��?%��r���S�T�� ~��/|��m3D&���,1��P�x�S�I�E�c�1;s����~9�?�ړ4�P�sgQ��
4sג��q�0k���;����=�	�� ������ ���۠��g����J�B	�J�T�+���R(ɦZB�n�����ً���t���������y�tv�|?G;��~�l�@��r�A��S�
�ԶO0ܫn�K��r���!M���N��x4��l^Lk�c�<ftb�5����mr5��AIg�z��1� 5~�ᖡE�$ 1����uF��\��p���_��w�w�i��2��5�6y�����ę?�dY橮��4����L�G�� �A�lچ�$wuE�Yn��Q��$�qP~l\��?h?Ӛ��@v>椒i,�h(�r�$7]6ؖ��',v8��s.n�]	[bi<SH�&�xO&�����|���v��Q�6P�^W���%�B������6����6oB�+�� �X:u����cэ��*+[�j�����ژ>�^E!��m��b�\!�7�]��˶�;S+��3̀���q*o�sm��De4�I�|�W�.Xk�D���{�vuB�f�n�S�;�ĞT�i��J�!��m�!�*m`,`	kQ�Ȧ��86�>:&��!�F�[��#��^F���:3�Uc����k�)"L2i���v��>�P�	F�۱u�|���\.����,[�����*_��/N����[xU_$�s��-9D:�g.���.n�L�6��(=OBF5��r]ޒEڭ�
���.��`Y%7��b��5W���6��Z��Q���0�R�I�k/�9Š*xɬ�D ;���	}�zI�9USW?�OA��!������t�)m����ib^ZƮ�e����7���|��0�q%�"V��7��XD>mY�E�c����LY���y�j=aǇ�J�;�e�?�f�U2a�m���o����<��D��=x(cB������q���P�@��װ�/3������٥�� �
��2������_
СG�k��!�5#���R���	���9n��,��Z�k�˒7k1�Cy�Uvo�����~u��zN[���;�Υ�Q�c;u�M�!ڡ޼��ɑ;zrݙVt�q���M�����g5:C�/��O�30�E��m��t{
I?Nྈ����,���
?&M6��cE�A
�Y�@�i�b��.�C��9���yz��p!�����K�����$�n�f�� ]2��F��a/d�<��
�83/*�d�yj�ь�q�8�lj�����Yh�����f�=]�=-o���N6�3�\�<�}_���n�Sz#����+_�:���$��ٌ?SĈ�	�]��L�U,C*����� �O�^ѽl[# :B�[ޢ����v7�ֿ"�EĈx��*�ݐV�פ�\9�B$I��6�i�R�r��=~3�1-����P���(��:v��'�>)p<�KɅƥu%'��6ت��	����rl;�W2i�+?II�a�X-�x�!��:hlK�����-�%7v,��m��9*[�u���_��Ͽ�~oT"�э�f6V ,ąR�pb���E��@���q��u��� �]��k�p���Z��n��_Ekn��K"�=:�����h��o�M�)�^s���\��tǹG�g�\�ķ���H1��������#�K�?���m,��
���Uݰ�&������tt���g�S��>���ь�u����r�ǳB�f&B�9�_���(L�J��>1>�1��gߑu8�]�U���	�E�7�q��w�ML-R���$��O=����ҰY#�T��P�`J�t3�i�Dԉշ>* 	wmԖɑ�C=�$8�]�����
ӓbJy���	�3���baԷQ
�2��-U_}����Z�
]���o��%�N�6���<d�s5� �_���ԕY,��{��8�>���E�l�y5����BL���_���$6��f0��l�E�$\��?T�&Qu�ʢ��Hb7���(x� �䝫�֪E��08<��R��FB��������gg�w�b$r]+��8�=@�J&A1�J�(��`�X6(��Ϻg�Q/�˟!�Yz����a�U@�*�f�����G�Ά�D�E^����dۄx�a4��Mʆx_�����bq,�c�)�q�Cs1*���
:�[�{Zo�y�~J2�O��)M9��7�}�SO,}۸�f/�r�i{KL�"��\߸[W���yy�r��MwB���s�&*Na|.=p�K��]U���s��n��y;�ʊ�׍��X��8���@a�@�_�!c��d-<� c�0��B�<�kb{�5GY��Fi_��TqU�'�
��MyE��T�˽�A��T슛t�i�NJư�����}%;\����\�-�ı1�=T��3CR�rqp���G* ��}ōo��(�`%J�9�7-QB�w����ME.� �~9�Q�+~O�=�Y�|S�����F{���z3w\��`dǜ����L�69������ [�:V��BYG��\w?�Vn����O��Q�_�T"υI�E�.�C�`��rHh�Y���ذ�7���+UY��wb~��òd���W�T�Ҿ{UR]=�(��5�KJ?dCK���M-�P�>�bL�E'0k�9XNZ�y*�_9��������;V!hh+;s	VVH��b�1&k
X�(���&j�d��CG�L����Z�Ȓ؇b2(SL2�w-�6w>���Q��3�\�8[�)c޵�2n�@��l�	l�FE�V	b�d:�~=��%ۢ���8��A�����&j2�&�����5��}g��՜�D3�>���3}�b�T$Bۜ/Tn�:����������)(t��I�<�U��0�8�!�[8g,�R�a����� ��X�c�&�V��s�c~Ȟm*eY�1��d+����������Ү�]nv�ݫ13�ު&Tv�1�op7M?�K����l�y��,�I�@�٧�m7��N�I�4���G�UG���"��"yyd4�l�(���R|���Ǔ�\���n����?
Q�1���M�>���"�o�1�b1j���!i���a_��0�b�!T�[U[�$��Ф���O��:q9E�DU"�-�9�q�p�\���~样�+0p$�.#.a��~tu�*��W�T�|�%l9h�U���'Xw���;���9-�^�k���+�l�`�d�>�
�{Gg����Ĵ��(����~����Z�^z��k|�
��@�c�{�,�!��� e͖9���W�)�xѿ��2z]v U��ab�s�I�5���[���˶��v��~@pb'��HĴ� t��w�h�3�E��LՃ�6K3��nu�%����@L��F{,��a�e2 ����Qmd����xiV�sy�[����ݤ���[�0�?9��Is�߅�Y75�A��p�E�>NXn�T��KV�6/XجVl���t7z�;�F.)�#B�NT�V����F=ʋ�I����v� �tR=�3��e?B������K�s"_r}�_T�"k_5�j�W���:zEh�'vC{B�]Pqd!ћ�%��+a�u�i(�|)I��Q|-A�Ox������8(�� �6������5���5���jJ�m7
��.0i�5�;�\��U���nnS#�%w���O>��a��9��R�C�
�� ˔քE ~�.�8�@[��o���/�~�ܳ0V0p�?�4r��د:=��]\��c"b�� +W�\�DD�?�ʮ���FýB[�e�'q[;���)�_�jKL/�;[o3^�(܏�2J�Dz��#�^7$��8�܃z sӕ������ap*����$<[�!��aJ�=뎩������I&+M�<BjC��u *{/����̐p��9a�l�W�Z@� ɚ�z��e5AF�2i�?�٣k��Xr�L�'m!�y>Nq��w���{���H�U��\k��>F%Y�}$Ԃt(/9q���g&�½��dT��)u�i$�:�xi�*�&E~pK�?:�R#�r��5��]�*a�b*���u���w�3 )��� M�
�B8���Q ~��cC����/5��� �&n~B��)���9�oa��1�*���F��rR�}J���Ȩ���F����aE�gy��'W�g|`�#�$ڍ�%��F&�BPo��g�Oy�w��c4��)��lw�=ؠ.�,�KH����T�c ��+����#�\�4Ǥ�U�K8�f5ٰ�B�?3�o?��dDG̮����`�Kz�ktƜ�a&�cz)8��#��ȶ5��� �9m��	�F��p��FC����9_�fΰ�⦷Q]�!ğ���O��N�k�;=��,�1�$!�V%�}K  �mk�=1%�n��+�)�ߖ����?�Mt�D&\����\N�x�^��@�����Z��^lQ83��1��L��6��%�ϱ����P�q�@��"@�b�C�Ë]�c�2��S_�W�:��!3*��z�_�	���G"�E�1� `���}���J:��r�/�V02��zb���v�u] ;ه|��D��`���vㅵ�������9
��g�g��_��v��Xdh+�B�AA�d+���o�ZY}�B�.���(F	=b%;d���E�g��!�,��[��2�@]6�i�ͼVV�������gyk�A�@-)�(��p=����X � �!�xV0!�Y`�����g^�o ~�����I�IХd�A�H�]��o���q.�ߙ��m�ilpG&�{)���"�D4*�:Kb�ܜlԉL fi%�������,/�K�y���%n� ��Dk��o�����b��eTS�L��4Ř�4uާl:��������n��?U%�8����)_����j�'s��Y�;�Ԣ�F��g����[��2bw��̗ /��%��;�)ZprR>Fb��d^ wM7�}y*��kX����,���7Ii �P���nFvn��Cs�P�)�>U$���K<�x8�� ]��(:�"[Ex�*"s,��׹XK[\�����3�pg��BF�G���R�b�[V��(�O�ag\;gO�	�ʪ���%2�'jܞ���6E��>�p�H��+�s� �X��5)D�X&��H��&�,{h'����?��Ud��Сܠ:�<KO�8MI� ��~��R��|F���4���FT��U٪)ʋ5;�����tJ��V�9,8dC_W����OY��&5fu�Ğ��@	��O��y�m�����<�Dϱ=�2'i,1����-l�L� �֠֨�MnibR��,�ɦ�pc?	���-��l'�ց�:�#�H�p&o]��.p�0�zO���5��g�[3��[_+��A:����	��ܮGR�y�G�)zķ�>����lNo�`^*dD���K�v���ڣ�9�|0^ʛn�
�8oR���=��]fu�ak���r?�5N
g�~!�@}!J?ş<��@�|�7t�	YҚ��b�,�Q�Z$3 ������xGyfF�{�B����������ڳ=cV٫db�Ah>����Y����',����j�]V����d�N{t�A��%��uC�D��my�Ys����"/4�M����ŘI�M��ߐ��6y�L��U�L�3�'�G�,���}����>_� �ͩ���?���pz�`��dG#v*4ͱ�nX�C#\y��e�ri����`�X"�ŭ��f��!���"�BPn�Y?#�X�F�����v
�q��<3 ��V�ܐ�(���մ#W�<v�ѹ"�s"_VR���;8�lW-FZo����
#���>M��{!�j�%z���E���Y�L�A�Y���8;@~"���i�nG�Tc#���z�Tf*Ы;Zot)73�K���Qg���x��|t��`o��:b2^s����R#MtE��R�yz�Wb�,K�sn�ȕE�K������~%~3�<AeL/FyA]�zd�D����gw����m�Yt$�Y�@���u��yA��)>~��bǯ�AEqc�{c�{upr8��r��.`y���<5��V.V����PԑP��?6�xUϛ�J�����EW���\y�S��?�	MU���L)�����A��l�*&�M�݈�ŉ@�q�K��7�u����p��5�-P�3����H��]���}xI�漋��U�*�~��H�5�����vol�)�3�>�S`�n�(���mW��L8��p��*�Y����M��7퇪��TI�Nc�[%��^Z�Ґ%~k�:���7��@I
9v��~���]��Δ��&+%�H��8|�"���1�j�[(x1ty#<� �eP�>Q�י��A���D=�����W�8��upJ�m}2�U�s]�.�����y��41�q�8cymi1U�V����0���D�r���@��X��8Z�7fB�� V��,��1�����#q�I��ܖX��J��	>��rGuR4nI�,H�m�mΉ�����qg��(�Ohcż��#Z�;���UL�Aݼ�$^���+��D9����.�Mi��]��J:=f4����Ms>Z�h�x"U��q����
|~���3l�Q�#\���7�'eaW��f؏hI��zI��j����ؑ��[d^�Wq�˥o+�k��D�~��uB4;?�%��.!2�A�yY��w}:�4EV�#^���D�sD�u�u��Z��ϣ"�u�9s���0
G.�"g��Y�1���f"E�k�v)�LT�¼��m�0+���!�,(� �,��uUv_.��{������m��^+�GÞK��W�%=`��`�r��y�a5�9�J�pz�֍2�G�B6�P
I�q_��5�c�����%	vg��ċ�l�m���\��Q�X�==��_w@�Vy2�|V}cbf�޹9��j�c�b�n�L�y�V0Q���%�a�dk������
l��ͭ��	!g���!F%t�$�#��|k�z�L�\�T0��� ��_,�9C���է}!�}�qQ�Q��r���#�4��� )^��{En�^��F�≼�癃�\�Ly�p��r*wI|B�E�ʢi��J�L8���L� B�AO��5��?a������?2�Xls_��#�5δ�n��p#�WG��F:��6������) {�%f)<��&�OE���=@E���?\������ɨ��}�!�}VV$._ ��m�/鞼S�$�!��Ett�ٞϱ�M�5�8ۡ�%;&�6��J� �L����'��4r��5����F=�G��ӵ��i|E4aӯ%�k6�x)��X֤�X��`�&\
䀪D�E�~�k�t}�KF�4)�%�ڻ�aN��m7Q�#R�;۟�%AZj�do �p�T���-V�ר��$P���j!�uk��H;n����JM��!�h^�i�bL�&0��	=�f�SfR̟�<�Ar��ÿ�f�6��$H��/%�/��h$�W9sHZ��lǡW�K��!��8P%;5=�H�wn9�+�fں���ة�z5'�J�')��������a$���&��*
���ڈ��b"�\;}1����;����������C�̽�t37�&W���Q��$�m��0��gF��Ç��fx�^��l������r�Jo��\WR���玽��p�����h]Ӡ�+Xҙ�[p	�:�'	\��vG[j��pi�Ie�2Y�_-��7o4�;��2���n�1�4�e���_*}V?@L0|��ͣq6�ǝ��il^E/�
���ǶME�1���.��:|M*3��ָ7�����@"�*��:T{@���o5�bh64&�Kջ��r�)�QD��|0���V�K��a�̸�B(�d����Ba�:�j�!y�����K��8Y)���Ǖl��A@�}*q�š�ɜ�H1w���t�b|��jj���J���#
O���Y/�����qp`<H1���y� ��-���`B �g.i�>�f�)�<�R2N�<�n�wx�˶]�o�0q�gHs�e����i��FYf�ܔ�3�v���t�R��<A;,���}w�aKU�ş]��:��\{�1E"�XՍ�6Z��\���{,CQ�-A�U��~YMJd�d�Q71�?g��B /w�y�E3���VW�z��b OlJ/έ�GA<P�y�{�ȧc��3y��m�KS��6��.�w�>[t1n��G�y�r����:v������#�hy͚zI�����-��ڍƜ�*�r���ÜS���8
��0�s'+�ʪY/�FBr$D��$��?t�lE>������M6�����Q؅��*�P�-��n�T͸0vH[_U�V�)!G�E�@^�[���ܽ�h�GLul�h^W1�����dL��f�/a'y�&��ES�}?,����(�md,VV�87Et r����l�rh�Vz_���fҐ���D_dGS�	��Ԩ�K|^Q�����o�Q��t�BC9f�%��;�;M{O��2��9n��_:#��m�1��I��".	 �q�����A\��~-#1ʑ��ܡ��9N��a�K��BϾ�NN�`aj�ǩԞ�mx�|�>4�/v���VA���/
,��Z�����UOЙ��_g->T-f�;K��(������Fpr����xM3ǸB!����)��F{Yෞ�|f����fLF���|A"<��� .����d��V��U.��b�Lb�P��?יl�$����be�g�Cp��z�Q���v���H�u�����	��)���i���΁��F��*��9�	p��od��L@�����!㳽��̙�,�BS��[��RY���!\�O���s��L���N�8$J��h�)5��|�r�U/�����U��L����:��`hY<�~#	��S�l�<�+�����I����J�u��%|nFؚy��<R:����x��f ���Xo�pL�9�����cE�2�/��	���%+��d!!��?W�pB>2�w�t8�N��4�p)�&wW�<�5��vvG�u� ��2N��Ĕ�ᤸ���~ ���Z��.�s1
��:�T1�Z�-ś󴁚J�ȋ�������\'�#g�s]��d;�I/��a/��A�ihaK0�q���������(�V0.�Kp .C|~�&����%�F��ƈ�������3P&��|j�-K6����.����zl���	���j[h7ۅR��N�:x���Kk�7��T��M��ێ�>WY����^*��jh��7`�*�l�ӯ��%҇9���e�����J����܎~�KV�(�[�}��"��`Q�x�j)O��������V�0X������p����2ͭo^pF�^�d����a��o����U`z���h��lKm|-N���$���r����x4��<��N�<�`Ou�,��[��|l��.OVq3V��!��������.�w'	� g��Po4���U�ZNc��A�ۗ���_m��b�˕#�5�irp��nMf6$7ƾ���<O���/@���|��l�����P�ߞ��H���k_<L��A�\O˴��a���Gso/_���X%�yq�2��vb��n����7����\lԬe�<�`:0��1tP�Q�}�Z6r�I{zhb����f��0�h�)O��6㑋-��c��dE�n���9!9�c�o�'Rd9]�,�xJ��yf�Y8`0��Ub�e~-��u$D�-д9%k~y�}�
�w&���@���~����ɴ=K��H�`>퉵U�A���v��� ���z�\o �|���O��Y��O"s������XE<���X�Fz�Xri����Dv�΢8Tw��q?t� �5i?`5��R���z�2��M�̰	bNgBJi�����TWg���0�Ӧ��λ�"C���r�ʒQ%ld��~�h׍[>\�#H�^k��t�{�PvMmsPK��4ox��*�*f< a;Y�Y�����!o�5zӁɎg�[�E���:�F8��Տ�dK�B�vr���+j�� ��KLω����B�8�ő�xVcj7h���S��L��`���s?�Y��hH�>�2$e�.uy��`rK�{e��?�X��
��W\��eZ5mVe8��f� c���������ziV�.BWқs60h�iOJNI�0�r[�!C����]��3=>����"��i��i�t&Hb�i��� �=s{׍�Qh;e5֜��1��d�B�:R=~�M4pqs}s��B�Qk\������ <j�׆��T�B�`J&rݙ�P��g7��!��2c�\Ӟ�k�+b.t|ì�^�����ƪ#:�/�N�����g�L/�a��C9	 aӻ�nt+X�ߋt�>�넎ȽSG�/��t�z�W�N���X<RA{G�A�f�Ӑ�8�1ۨnKt����a?\نBGv�/.ƃs@�<���XE���H9�t,�깎.Q}���� |m�ӎH���x)�Z��D*;b"
�X�W;�S�����.�9I~���6?U:!�6��L�^�[~A���Z�;������u�v�Eawp;.��n����_�#������b�u��h�,���m���x�7V�^)�E�z�_"�b��s�f���C�2cz҆T
Xnw���9�h�e�����b��T[Ȣ����\�CU��ܰ!��6
[��UF%�����>,t!���4q릍f�i9cޛo���{ԣ�?u{x�;`4���jT�ZCgo����L��F�?��ϗ�IgnaR��Qf�73*21q^M,��v���?,�Pܠ(��F�y=�O&Vm���He,T���gMg$,%T+��z$�]I �����o��#��q�����e�-1 ڃ�A����O�ֽl�¦6jG뷞�c��<)u���zK��WL���=��4����Typb�
�{��ޗ:�VL��m<@�;�)5�>(2��۝�� �ƯđN�-�ō������U�֕��S���8����.��p-�,qn���W�*����R�t0z�d�C��T�h�&]F	��y���$��}�(>k������εoۈ�Qt{�/sr7T�,a)�nW
�8
2>;=Jsť�	G�g\�X��g�7��dg8d
%�}�܅@2�T5#��K|؝UD(�k�~&�
x�����y���M���s����LR�/�c�{��&�(!�oĆ�����[@C'r=c�P���j�����b��[,���z�����>h��\z	�g�M�R;�5�n14/|�+�����\��M��ʚ��ꋮ�d[SQѣί6�P
��3��R1��D3��� ;�� �Z����=vi��H̃x�.h����K���:�dc.<�In��z��-uA���Y֪���b%�����[.���ñ��fK��O�T����u���t��x����K�I>�,&N�A#D�H��P�����;<�P|�)}O�T�0�F��F+Ǭt.�oI��$��/^HgQA�5��re�4���<R��B��ɴ���	j��v�4�/Ң �c<�X���"V����l��׶����
��%�dԝ	�]Je�S��5p�`�Z-��2���v���&���zx^d^;2���;=�!+$�l�<e�E1�|����oН�CHlBcv���&Ԫ��괝
'7��g�|P���Qa���� ��f�P �h�@�A�rڎ��!�O$]д���%}�޽u��ɇ�Ԕ)ȕ��o"����cۤ���@;z����n�~r\jO�03:I2���<�V'�, 1���Ei
.�y����iL�c��:7�X�����>Ē�B���i�n'Iv��_/PT51��:$���َBH�J��ql������˄4}�H��C+ˋ�I���l��v�s�:,b=�u��7�I�����@Aa���=�z,8�S"�q汯k���U�9��&Ã�lh���һF��C�%\���3GRq���ۤ);�۶bЛ���0a%S�h��������0-�ԍ���E���fy��(v��.�Heםe��R�3�����Gj�Κ�^�p*Š�����pb�^j��ȄF0V{�cj@�b�����'OP��(����S=�;ρ��:�h�թQ'��O����+��na�A�q��59�ʨ�Lk�{]]ʋ�B�
����62�e������<��yO�Jk���f��b�g�	m��)�u��4�3~i,[�[:�F���,����S~Ӯ,��]�y�t�ˢ+�z���զm_/�D���u�>D���!d3������|6Gy���:�!��JawH�y������S/>ќ��6*\�a/��-jB���1��8�U����a7R�,`O���u�$�����ŉ��-5)�XG��jS�3�;�Əz����퇤́����j�喝��(@�d6e��=� V�pӴ�lL7��bed"/'ܨ۬�RF�m`�� ��㋠����������U��~w��d���,�6	��A���Ny���:t
Nq]^���s���}�,hפ�g�Z�fjE������ܙXR;<��g���t�Cҏ#8!uA>��s��a�ܧ7�#GY){~RM��8�����ҳP�m�eb���p�5�r~�\V�4�#���¼.,��'� �We���@�Y:�U�*H��:��.��b�>(�;��X%G�LŶU*�����:�����`A���4u�<E{�p[a�q4"C8��g�^b|���!s��{npN#����٘��`�6<�AP����m�X6�};�,��㠾޺�k:S�A�GB�%���Ŧ�ByY��[���)�Uj^�圜^)��|i0���m	v�/�Z	B���[�o2��&�ʊS}M�R���I���}T��M����Ho�\T���0\%�p�ߞҁ��2y1꿚g�o���a7���8�9A���\�3�0�}������Dw��5�=E��.�ڤw��A�鉄N�<�湤/ێT�2ު2�(�eh��Q�V�	��m'����.���6���� �.̷��ua�u��@�eqDy&X튀2|��K�kO�1�-m���,�=UD*�0�V�x�>"��W���r~����tU�6��Ыl�/"6VM���o�N?W�@�p���~���1S3V����v.�F)10GhS�-+M��_0Nوu��@��∼��U���Ʋc��N�����;�tyI��&��_�&_�t�-�v�P��9kQ?��en���P���1�jX�K@To��2Wec�o��>��:7DdR��L%��\��z��N�^�R��h�g�������)�ڄ�)[�����>���w$a�OR�SxҏA��{�� -��+�3�0X�a\�+��ֺ�;D�^4��᎓�z���T-�F[�����]1ЍA�k��S���3\��t�o4��&������1�����E�ܲ�_�s�.KfO���mPҐ���
��rߕ����i0�i�5H��!g��}�P���0������Ɯ�6�OWʭ�;�޾ƗX�l�����co�&�QX�[��r�2�QK��qB�'�t`��0˘�]�����|+:��k�NǑ��]{��pɝB���[-��g�)9uzD�}�#�f���o%(�ɹ�
������xO$��+t��8~&X=�p�vm{+�#��;��lX�l�ב�ٖl
�O]���f"h&ڃ�0[���8��7���(Th�n>]F(|ڜ�4Λ�+k�J���R~2]� ����jkH5��E���E)Ҁ�u�ƿ�a^�4#�Q5�Q7�9��A'ԣ5'���:��rk@�����pwXia^�Bp�;�}|n���x�x�c^ �k�:�j���6��_����*��J��壜��j��*��/��gfi>u�zk�V\u�嶌�+�t�	H}������.õ���g$ߣłQ�y'��I��9����b�����1F�npE���KpU���jh��;d����~�5�~�8Y��r����M'��N��"��H��N���������������/c�ב��Ӥ�뗅�N�>������w����=)��@����z@r�e�\�[�gsj�l�\��'��+�@���#�?P��<H�O�F�.��.��A 4���)�V���1�}#9����%����'��V0Mj�c���V_���l1���$���q��fТ�k�H6��:���M�*<�[�����bފXa��o'Tn�*���}����OƉ��kA��/N�VX��߷�y���j����V7�I���� 
ȱ�_V�%�p	��Cz�q{Zc�&��v�Bls�|eǆ]���k�?�����]n�B�^&kε�L��f�����{������9�>��N���t�h�cQ�3��/G�o�Sa\��çJ-%G+Ɂ��&i��+��b�}��,�7��0��3� 
����k�)ۛ���$םA��\���[Cu��}��\jh�I��R/w�Q	*u�A�q����L/A����@���kQ*R
��bV+�-]�$"u{�FsC�A� �ԫ9e=)bE;�L���I娗�2�۟1��}朿�f��ޛ��V�c#j޶��hAD�4`�׷(I�!�v�9	s4��{eؤ,��F�V�W\�S	��Ȭ��-��[k�y�8>� �(B<��e!dD�p��?~��g�:�7�f+ b��x�A�3��h9�,��>�"4]�g$4ijy�v�v)��ɮQ���?�I#�