��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��D��ÊC�f�^����mq���U�����f�>�~��i���W/����+��b=G@\�D���>���sL�̢Vh��eP��*����v��Q�D �������#;[dM�`�����<PG��&��l��H�Ɠ�Q�� L��6��I�Qa�a ����N����*���n�h~G^;�QW������������?G� nE�92e%�t���n���x�h*�߉BN�p?ma�(�zu;gf�.�y�>qv��b$u��b���F�2_4��X=�~z��=�WƄ����N�[��W��5 H�?�=(~NՆ��:Z�UB#	��.%��>W��S�ĘZy��Gu��?J�9�y�	d����uU��5.��������6/-B��&_����� FM�S�2��uS5�xO,��/�x�WOi8I,r��=#?�d��y[f���,yB���lP����4*�6X5\ut���Jca�ޙ���tO��1�_���m�0�Uxnf��0Mԧ}0:�\��$J�����͕�,��u��Z�?K��6	�����5<9L�9D��=�?>��OD]fTd¶$t��+��ovH�N�$�|���n-�dp�V�ɾ�d�8��������rE�x��^g�&��,�����O�jcP�AJG�.m -ބX��b&KkK���j��m�n�[ĩTÔ���r���%/�{��a!?�T�<���Gets«�Ě�O��d�w,��ă����ſD�2GGSi�es�G�3%(�
*zL����y3ձC���1�OOD�N�I`�F��M�͂_��N��ϋ�8�2H��4/K��j��b��w����A{%����y��aF ��2g���g�cٍ�M�>���lj��4c=��H����h�S���E`��e���,}y�:iC|ZI`yT�R��^�YpF7Z��+^�
��8�~���Ȱ,(	���a<�=u��i�<�xi aoޥcd��X�I�K�r3� ]���C���
��ګ��z�9�۶��F�|#1�c�š�{ ,��0�D�Fu�I���\A�2�����ɋ�D�牡x���E&T����v8�A�6>�5F5!i���}����q���;X8�,w"�$�����.45��/{�jP�(Z&���b���{
�.���VQ�`��Zp��
u�5�Ɏ>k��~�j$�2���}ZMнp�jŠ�y���-�襀S�r�����PYu}�wk�a�ɸ�}o`Cn��Lf�n�᜸���L<���nD +ޭߌ,��,���t����q�퉸��l��������k3K�bѪx˴���)�3�b0��\���F#;�E��F9�_uYi�B���L�5d$�	���I����aݵ.p�>F�ad9�ْcF� 2�YIӴ���	�+|�X,�ޱ�F��l�D����2MHUs���"��7�ҕ��h����T>c�i��ўz�2p��'��M`�	�[](�PM�Ut��V��Q(�,�k���[&&.�L!3�Y��-c#=�]��B�$K,�%K�h���\�R�����ʐU����r��l��I0.�����,���O�$H_^@L�n�XV�ʵ����ѫ8��wӯ�l;i��b�q|F��l�%W��y��������3:��ﮅ���󎑻��?w;�Bg6���G�DӈՈ#"����tO�p��0���<}�#��-��D0ֆ<���TΞ������`�����莏�S�q��H�w5�e�u�hlo��v�!$�"���#�-�섀
�)��r�K"Q�F�?`�����O�\p�s�r��a%�ؒ�(����M=�4ȿ!g_\��K�$E���7f��Z�O��6<�����Z&Y'z�B�G �T��0`P�/�8B�o�G�RUͩ,*D�͈2S��>�H���\��Q���0G�����ʛ���x�[�#���{Ab�uG(��k��h<˚?}4���u����V��q��;�'Ǚ��T�aH:v�D~�a��ە�!U��'����O_�����*`���`�+=�gj����r��=y�q`���!C +�5�tm���$U��h��$�;��G̓f�l��U���N��.p.$4�n�@A�sq�kϐe����$Ӯ�$*�~�-�9Pz����kD���i��,r��	��w�bx��b	&����~�O_�$�8�#A����#�M)C_J���I!rcb&�������ۧk,8��^��1�!>�E-������N���3�K�`E�R̶6�����ܥ�#�~U곁�P1�e&b��%��b�5J�<Sk�aХ/��~�������z��z���MB���!\��.�^��`j�ePt�5�@!w�XMֳP��X��� `5��Z��.�w�7��B�C1tDs)¼xD>~�B����^���MY$c�5=O^�oeq�lI
x?�C5t���L���w���&SN�%_,	�F��'6t�����Ww�i#�l;$�ªf���53�
�*�͜C�L�s���=��\���1<,�+�B��.�/�yMf41�"��}�T����`�q��Q�6i�����۹˞ظ�٭J�`[���w$K�����X3g��Z��`u���z���<EG�L��k){0���:E�C����$��Bo����d^��)����՗Q�m�}�>X +��mS�e"�F���S�F\�qnS��싎��
M��]�M�����������8y�B�A��L̬K��{��e pl�?XP�#h���C��?�b���n��j�$2a��7���͔�c̨M�B-�JG�:��h~�C�,ĕr�l/ڴ�p���xO���T�k��C��7u����*��l|�EDm�+��Y.^g�[���k�=�	v2ɟ�uʌE�-�w�	XD��ޫ���J���0zoُ+���US���`�E=��M�9TÈ�|��(��>-��P���v&,�L��se�Ɇo����� �w׶�isA�y�F��<�g+H��o"�CE�n:w�de�5�>L�ͨO)C�T2�뀨~����~�}���^���x2��CO%/}��(cj����0'8$;���~����!�QO�.	� >�f��Q��HbGܰ�R�00�Ε��7�}n����J�Ms6�d�W������a�,��(�8����ٿ��ط���{�J��s��̏�R�'ʹ�V�~s����6)5sK:1�J�B���n:6K*7`B'	;ڞg�����[�9��� kLM�|�G)����҇l��OAl��mN�#4�ژM��C�2�}~�Z��cfq$����dc��)��'��e>Y�f�Y[����	h�j��/\�p�h�<&�����C���J�$0�R+�]p��"��=�"kd_��M���tQ�;g�|Ma�o�b�Z���_o�R+]��L���MzL��PBY$�q�G���n-��!9��{K$�ӎ�#-�{��&�:N]#*&�PCm�$�r���z{͏7%Q@� w{�Y}��W�ɝ��U�[�Zʖ�%��#>���������9���ώL*����g�H��4�}��ғ��%6���b+À!#uJ�#Q�-N�(�B�mq���I�19o�Ђ:c�����Ŀ����Opr�U�l��X4�L�D_h��2�	*YHǰUV>9����K<��g4M���A,F�����S7˜N���1MXF0.���\3ʯXq��v�đ|��P�۱��I���,u�K�I�^��f?�*K楕	d�8)��CI ����z*=@�U�}Z���Z+�K[1Q��2���~�+���(�?����}�v�ә{x�>��qi^�H��A��Nb�0j�؏�ye6�7���η�kY	]z�I/�g��kH�ũk�-[�=@��r�[�L KN6->T��X�԰�2�x����媛�@:��|SK�Xě,,
� /_��t�=�����z��c&��N�s=��YeS#=㩞Tj{V��N�;���/Vt�N���7gh��o$��F��M�6��<���ቤ���.j10珑����I��9R1����8����|���|'��9y�x��Ë�����+�F�`i�Z<�Y�5v�ւ����NW�:f�WW�	�++��vR��|�_�^�ýc�A�;D�����_*���!ЮH�������&|�Ue�k>tz����~�/���k��ꚋ`������7�:U��ݠ�"s��I��;շ����.:����Q,�=�x������Z8FMgZ���;��:����D���uL������v�H礧ޙ�4��)d�G��4kF�Aq44b�����Q�f��YB�����ھɤ�,qq�6�I,�T���ڣ���E���'�~G��,�ȫ��#V�r���)��Qy��|�|���_i����x����E�)�%��̹6��s%�Ȋ"e��wԟ?�1�3zqm$��/�|�3˳0�@?��7X����s{Ksh�ؚ�����>�?�ΦsW~��h+��uRR���2���5���nm�o����ՙ8�8���Y�g���t�޴UQ�X�i|wߛ<>�ڍ�Ҹ?��N	\\=�IP����/ղÝ��]��"��߷�	jW��$MniD���^U�R��,��쾌k��=��7�.�^5�W}��c�O������t~����:�?�,#�uXkT��}滮�'JD\����vb�3)���J�F���c��G���(���n���Xկ�_N��F[��c����N�I�b�ݹ�g#��I�앟U��m�-�L/��rw��6�Ǝjg �t�%PMX+��#݄�:�k�޽y�J r���`F��jwj#�n�帊�m�_�Q�Ka����z����0����M�	P�;�Վ罟�Q��}j���SD�EY�%���4P�Y��e�*V�Ԫ�,�uM�Ԓ�:�K��3c�f�����ݚq۠�t���K4�_�^|�q�L�˧}"���f��(����X���m>~⽀i��(͟��}�j�yvw�]�,��x� Oh�by��gY��Z���̩#thVX�鑚������U@Ι0�r���1�x�U�Ѽ��K
ӛ9_�z)�����>ck>���@�j �&D!�^�Q��KE5r�S�7��˛�:I��.r'
2�7h�X *�
������u��p9�N�Ն)��'K[Ԩ�#�_P�
������(	�l����h�R����$򕰐{�p�;�BYF��7|d��F��/�G�"y^�4$�?��P��h��ƅn�3��33Y"P���Υ�Ύȼ�g����$sg��Ֆ�xa��i���F��[(�%T����+�]�\���0��#��y
�1_��pf�n�B���
�Vj�B��y��4�uk�g5i�/��H��X�T���_	Id��e(�~�^ �W,}�C����.DU�8�l 4��ii���9D��+�Y�
�x�g}`k�֑�J���FY�7/M��NC���U\��3�����L�v���VO��f�l��F��/�*R)�̻�����`�P_���A�o�
�:���X�k'd��y�=����`��]I7a�5U]���`py��ӡI�Q+�{��#�(Wd!�Z��?�N&��è���l�FL4��(;�q��,ڊ��z����c/�^ۘ}'�)YWG4X0�#�F�Fqs����O��m�϶�.�j���hcW�$���R���T$��j�P�_�g_=6��>�`���$��x@we��[Q���q�	�[����%ϸ���$_W�ZH�d��5r�\�D�� �7���km-���P���2.ʔ}ٞ�X�"���M�J�B�`=�l<��$j'x�A�Z�6�M�vk�O��i4� �B�/���)ʔM(E���E7E^tV���;U3���E��W
o����@������<�o�{Od_-1]Hd�3;������<I��=�y'D�����X���w,�4��jefR(�W�sd<��G��_�'�_X4k����톤�����:��*���<�̻��`�6h,.�m�lV�X��I���K�$���mת�h�&�0��v�(��_@��hOJć>�>��&&�ht�����W�:e�*�.�.�Q;~L읣�&��Dp�O�f '�>�������+T\�791��RZe�K�u�	HN�-�i-v�5:���b.U.Q�y����n=C�g����uҎG�qm&Y+�e8��9\S��n��l5�0��Ӿ B�&Õ�ەvf�*�PVI@g�)c���=I��*KX���,^%�	Bf/��R��
X�4�������R�݈�������)a�9��K��F}��Lbp��>�]�M�l�w�����HL����'Y�w�\�t��7?�y\oI��l�.��0�	��5��A�,Ye�+G�8/V=D�z�x���Bf�/ˎ¢�+�/�I��H8����E�����4��۽e�H�C�߬�ǆ�gY��)&2O�L��ˍ�8e�U:@
��dcT�%��9���,�q�Q��c4RH�iM�H�ۭd;2*�y2��F70�WUBp������].]�C����={���:�G��@��Ӗ��{��˽���|%o��aLy3���,o��Ů�$��:�?���[6�������r���c��T��ݺ]yo�"�|� �s����������(���������-�n��t7�|�8����[�4���M/"J�A��<���2'	�t�`O� ���	}������"5Z��(���\��s�{I��Ғ��%��[7�`8��v#@	�ԛ��I��v;"c#�#��%Q(UA\��2���h����\/�(јu
��D�^#�akGS��O����0E�xK�
�2��-+�~��ymh^�'zH&�%�����W_���D�OU� �L 3��,��>.�'�.?lu�Ań0J�<s~!������oWt�,��DML[���b?�h_��F@N�]���6ܭ�sSs��L�w�e��a�"��0[}�@v�v�E���"8�)�m�f�%��v�wz�����)���>�f�|�sT�Ϣ;�h�_��Ϣ$��J~qv�/�]��&,�M��)� ɤ��! ��1�?�1�U��	
z�Q��RP�8Jn;O���Җ�����lױ@�G�[&�__������ &��Z����MZ�ƶ[o�c+������X$]n�b���W�y�y�}��4��<0�h��1�}�AR+D��I6[B�k�*�'n�,t��
�S��$���VD��ߛ !�ӿ�'HR��#@L�L^
�9��#����J�v>dјPL�%D\R��9JjЌ�P�_�ܕ��H]�I�zU}���Z�󅦐��KC�*���;=�-�fTd�J9w�+�)�@��j+Y�t�V	sʠ�vj"z�faZs#�J;�O�AMEh���nF�]��!	y�m�yʭ�ZG�7h�2o�n�{F$u�:��/�4'5S_���k�ŎC��1�Vz�6��<K��J��BI9v{���#�Giy�>W7Rh��;j	|/�xhUZeP:] �o;����@���5�fGSR�7vef"X�t%O��B�߮%�,��yH;�,�zj'�����Qu%�f~�j�%vj|�pke� ��$]�fh������_.?�:ҋ8�v�Sw;�Ge�{T����'I��d�9�@B�V�p2��P��Oc�7�'���]�i+�(�q�K�19���|_�F
Qf�T)�W�O��ɴߧ	k����r1e�/�n�T_�8��#
�_�/����Z�*[yL�p��>&�W����>�1)���@�"��;jY+��'��R�ϥ�\G�@�޳��uN�