��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���!<So���2��E�!�7���feI�R�34�F�\1uR�XO.P㤳��"����(W�����Y�us�'�V6g{���/�Y�^( ���Ne�[�����8�1��{SZ�k�eZɇ�FUHn�i!�kO����r�o�40e�@�̺Na|�g|�O̲s����_�oW�h+c�	��x�1C5�]�`��P�#�Ι��;<��C������^c�4�\us	���S���x�~T-���]D�lK�c/[G(+ف���j�H�3!`��|�V�k�)j���Rrj������+!�m�iS�\�,�D nP>�:V0�(�9��O�Y����m���7Ӧ�J�Ā7��-�o�6���d��iP�2I��5����^��1֐쬳پLƑB?�(�x����wj�j[p��ب�Q��8�)���b' �{b����Z�مIt<8�3�\;++�Ҭ���7���$5�?��Hf���*"��6u�Ea1�Q�g=�f	����%'(�l6���g�L�YG9�:x}�� ?d,2+5���1;T��U��Kڐ՛vN��~ō능���d�>��$�s�D�Kb��{��V�L����+��6pM�ld���v�0f3���w�ہ�V����W��� TB�Ov�4T��9k�m����Ҟ[Cṕ�Q,:/I�ff7M�d�$#*�=չ/Ȋ?@O����-�+�g`��0�E�΢f�Ր�#��l9LBi�-�.�{��޼W��������Jx�a�8T�r���ŲG��@�.�f!`¾F��^~�G|�v �FLN�j#!Mʤi��ɘ��R�������L�"��[�V:�(V�R�Н7�i&O��Q3��������>ac-k�cq�"B3Вa���-D��+�;�IYd�xޱ�T��F�A��Ji	���π�[�>pE�����ðh7�A�P5�f7������:��_m��\󔊁��?<���5|���b�P$1u� �,�U�����Q�	$��/s�QC��Tb�����nO���n�E.�|�@��}�"�^_"~B��F͵�U
�Zյ'��^L18ik?p�:�yo�K���&Q�V��b�՞�	�Ja�2��ň3�����c�R����k���+�T���0����=A���6R�3��V�$�&�zҼ >m��L�3a���rL�hl��;3U�Q��da�����"}�47`T���פ�����=;fg�b��Z3���Q�-�Լ\��ߊ�;a���$��I���L�K�.�*i��C����wәֺ���ux��cO�L�xE�ҵ�ad�V ��^��� ��(���~��q�����%c�̥H!d���%��z��N�S]ΐW&PH�$"CDbd"��HYTw$���P�#|��}k~o�/V�S!a��D�r�8�(7+���"�ҩ�2��iWRt&�E�7��I2^��%�bK8�!f�-�7��70ra���v��� g^�(Bx��#��zi��愢�X����X �v���vW�g�r$R9n�r��Z�,�aPŅS��c��nrT��D��U/<S�=�ىI��<�GX:��<�H& k�Y���Tq�4Klx�������
ׅh?yA ��P��J�yX�Y�>Wt�,��u�?����e#�>� �E��!&���<���ܘ��2����~�!��HD��zG�w�ܸ�׸6��ݱx��j.L*����K-�@53w�x�j#��i�Ӑ�j;`�9�W|�wn)�>4Cu��A�ˊ���bnzo����\��,W�,�D{@%�7[@��4����@�B��c�dN
��Tw�ؑF�hZ�J8�u��6����8��@RF<cB�K?+U����=49����=əY׎V�\o!\WEK��
�B}矻q 5|�Fd#FNQ`�0t�`?:��$!���R�R���Ar���o�¿�s0��L�������z�3%}���9�o�u�!S��ޞI��C_��6H���/�}t�0'���V��ʽ���<p�+�8��o�ʃ ��z����!?��"O�5�Ŗ�(c�{.�K�K�f�`:`QM�Ѻ���2�� с1(ZP��f��(���W�����������a*�#U��*�߃�/�o�Sd��q� ��x�v �� 1�7UPrO$��g��v�FӔ1:nŪ�0a�F��*����Mj�9c Y��`�z`7p(3�H.���^M�>\�FiLj�J�(E{�fr���#H������d���Hr�.�8d;kT�T��N�b�����������?D�s���L� �
gn��;���C�p+%��4�qغGT�R���B��y|���>����������#�.�΁=w�4E����=ﻰ>��_��{A�[Y�7��F5#ƾ�OpK��F�?���H�i|���VO^W�������H�ӝC?�J�v�k/x��=�#I�hw��J�̵�7�ioi��$�!�H0#��#'�U��̓���t�5��՚DÞQ3�[�I�c��7��T��u��V��Y���h��{�#����d��@)9'�G����Kj�D��n��q/�k�''r�K�����MR�;���uЪ�Ą2HyD��12��ө�^C-���U�v���+G1�~�6T�L;Ma,���pG�7T���ҫ���������fX���K���#�C�o~D�JnD��Y'B]lmg����ǧ��vQ�WY�R쬽krm�qn1���S&�� �hi���Z��*��1�Ep([G�Bb"�ֶ�ǁ8!0qM�Q)X����\�5Df�\�W��gF����i�;������Mz�G{���C��^�J�u �=�q���Q��y|�pfv^P$��0��W��,l�>����W�U��VIa�� �gi��{����{OT�-H �QdM4�~Z�]
��T�f�qO}R�'搘8���P&��Goэ7����Z�1H}�e|5�3��t-���fAu�3t�O���6F�-g�T3��� $�*n)�����OvtT�*��:�Miݵ�{�gFX\��q.LFK�ʍ
 �>���t?����!�=�����P��jn�!WA��ݯ�Cl��L!���&_�@����N"�� 6Ux�h��8Ab<���%�Ai��������Ҹ&�|J�Q!�АldUTa�A����z DG��Y�Z�)��X�g8
�����Di��MK=PFF ��Y���j3�O������6���{�Ĵ��"Rm������G��DN16{j~n�1��E�Xx�C$
������<�{�����:1Rt!E�*u�M�@����K����/��l�:�0�6	�$�l���4��l��?��%pܓk�2\r,��U׸�)H)�Q��H���˟?�O��F�0D��o����i&�$N���X'|��}��$9v�|)ٖ!���.[�خ�\gQ1�$-=��@���@�MFj\4c+U���j"G�}ظx/�����"'�c�%3�Lb1��1�N|�z��Oj��9Ap�ڡ�Uo�~�R��J�f��X��i}�P����d��B�/�xBQ��;
�nj�_�{��(P�
4���5�!},1�����hy��cQ�ې2k���0[��*X:>��x$���"����,����t�H�==�������]/Z4u־sI���M�,doK�.��2?�G����z�$����b��R�knx�"�6�z'��]�P�ܥ@-8�3���S�&_AQas�qڻ��� �b{]��E,t?��)���|�vt�R}9�S�s@V5+@��*ycY�
��윒��u�]�����O�A�lͿg���֧]�E��r���I�21	�<�C�~�A���o'm2��Ҍ;,�MdZ�/o/�r%� �X�v'��Q��6 31��V��gg��g�9�
��1�w��$��6ѽ�忦��2�r�M���䔰LgZ�o��d��F)�^�=�L&%L|�Y۽�����XpLp\�5�IY�����m_z�idD�-\k�Kc�޻�^l;�C���Gf������ ��7��G��؎�nve�ܗ��VP����8NN�=)����JJU�*1�=9�J�,ދ�Yh���{dp��'N�
��_�%��fO�zM��<�����٠L,���f*��v���G9��$�C�^,�>�o[�,�	4(�	���
g����>����@ʡ?BzoOa�Q����:||L�!~����״o�[=OeAl��G>*����뷁��2��:A�������"&��9Z���Ob���wH*���
R̯A�^�R"�s�p�v�]��>�/#қB���\��u��l��'�?!��!]�Nsl𻢜`V�m�KD9K%�؃`����"�8̪�ޙ���d��{\n������?�(�i�_���EZ�sCi{af.�ڌ5�_�5�������Y��(]{4��u�}YN�U��;�#�h�-�.� ����/�Pmoj���(L�W}���N���"�&{��M�q�7r�.�Z#���nJl�
��TX�ף�V�ǤQ���ON;-&d	W�Ƀ9���{	EGS�˔'*&�����G��.�G��9����M �/��ʤ~LSJu,��0��"L���{H�.��`i�H�6	0b㲙�ڔ.����uQ�ߪ���%g�F�)��u��(ҷ,��_p�l�O��2��B�~�˿�քh�b ����k�S���:��L��9J��x'iA�����5ӍT����% ��]&��P����xjC:sg.�4�쫩 ��H7q{��:ϽY��b���!�=�XXc���2Ű�*�ɧT۫#���L�1���SJl��8�Z6���*_�x������]�}�uJ#���te ��nkt�'h��
[�$����R��A�k���>?��ux�TuveίԕՁ����U%:U��ҝ�v+�@V�mh7��_��
ى����0��49}�n���G� eq9YxL{p�����^~��X�U�aOǝ� ��?�����IR0���)ՙ�fӕ���
��%��龢������L�i�EūII�u������+�b/����T����E�э�\��v��2-��<�\�|6���ޟ��Ll�¨�-*<���U��(�Q��@�|Ћ%XQ6��k�aO��CŌ_�"�E��g2z�o�pxB�ң|�KB�q����>c�7<:
�m\�>Ji����e��x�#]^�cBS����v��2����
��ON#$�9�_C�O����*s��J�Iw�2��C�  ��*��Z@�������_h���+��ҥ�F#��ӎ���1�W�(;�-�x���ƭ;��`Wl��@��[��=�F�o��5��e\�C\(s�6��(H�=�	QsG��W����F��Y��ѳv��.��)a�]c�P�������P�a|�a�聵�zj)-�[:�HL��oW�n.�z�`Hd5�hs�aQ���{`఍��U�:�����8�� ��:X$����>$6^8NU�Α4��j��E����:I�?������V5���qi�{{7^���s@�e���6�����,�Ry÷�M�h�cj����<=o�R���<9M�X�5�Ml� ��� ZbH � ���活�у0�|6���ް�3M�� ��L�Z�ʘ�G}��4���޵���?�Q����5ęx�-8�ÔY���̥����([��'���H%���T6��Z}��+NLW���h�)P ���a滌m���c��5�~��N��]f��8����pT����{k�����d\]ԡdb�����L<���΃N
��� <7�6M�d`�2���/J6����,XU�;�ە�u�5�����Ǌ�����)?��"�P#,���fv�2��"�c�$��/h��.@@;��������M�����*��j���������-{m[��T���yY�2��
�⍁Tsy�l� �����/�D6��ԿB�Et�@4�֛>�v�2 Y�X�W_�ۆJWi�0]��G8_�:r��V���̔[�x���j>��c�ୄPQT�_�����4�C�,��Z���P�2*j �I������Ը�ep��r�4M%��1,��PEMH�S�g��`�Zĭ]9�ǐ��u�G����O��T!\s��Rrʛ�/��R�hMY����p�5�;g�Oچ�&�D�m3�<�gWmd�0��f���
<42��pζE>��%�K\��
N�V���}D��(���H�> ����YK����0��f>�@��Nt�E�X��~LM[՟3�ή�Yw�б=%C�/*X�u�#�ebA��p�QD¿=��C�}lA3��J�i߁�A���_5��p��ǁ��vj &����l%=O/������(<��ۅ{�DYx1���g�`��Ն��sIo��,�'����i_F�^9z��t� �WP���Xj;��ܢ*�6W�%S*�ǦZe���&>�QI'b	��Lyެ���@��[W�?��)s�A�g�8��p �hu�r���X�c��O]e�t/�W[؎�-�''ƌV���!��)!9��T���%HbM3�'�<W��)��>��F�|9��UJ�4��T�VJ�g��l�/Y���cv��B�Iv}·v�o�+.��r����1�A{�.����Q=[?o<����CO�J֗o�F�TCB�wGt�ku����6��ϕ�G){��-��i�V�G��OG�,,�B�rP��:|b��+�.~��+��8���0>`F��RH��/��.�L���	�!r�?<{m�ۢ����JWY����_���N�k` ""
����-�������G%���$�N�Ƽ�,�E�h�>W{��2�h��;�M���5�a]�.��PQ���R�L�y��X�"͍�+�/=	)�	d�z����Bl��c* �(�.sS��->������0]�/4�ZV@������bv�S�7��2�%����c~z�c��q�EӦ\
9�W�@��A���;Eno����A
�H��(%�-h�;�wW]p��CZ�QQ���>̐}�`#����Q� �Cn�vW�o�����	ʾ^ճ$�p⪁��w�OOpm��Mk)��{T������e�c��Հ��㜙��[]�a��i���2��/��N�h��p�6�	�	ج��X� )VI����+�c0a�d�����-������
j%�����o�$1@ i���;�Q�?�J��@r$�l72t��l�ߡ��(|K�߄H�Xc_��i�`F�Ә�h�a�.RO%`O���pf�n�Rs�~!O"l�����ׂ��2׀D�Ȏ?eP����K��a<��RVO�W������-vq�h`hT��F�􀶕M�Qlunu�&@��Z�;OZ�FA/#�8�X�3]�0��\T�{���7~���j����?r[�Ӆ	M�^Z�������y����W��k/��4%է&�d�D�Ol�Yo�R���k��]CgL�:x��Q�+�=dw��p�_;������A���1Q8 ���Zy���ӕ8B��dʺZ�h�Hݝ�ا'���x�s�G_��~:��R���qf�����)q��8�=�X���.�{[7���!.��&f���f^��",��H^�t@�[��SHm��ߩhG!��TSy�Wۊ�j��+��r�������5�],QoZ��?�w�\8�J7�;��?���-�w�T��J���� 9�����c-�4Z�Zl~!�=� �v:�8J�
�"`��E��"��>YWޏ*��w3��Z�6�b�ޔvC���}N_O��� ˁ�>nHfr�T�Zd51ɐ��OF�'�,��f�;��8=>DzKXȂ�7��_S�k#7�f�~�AXX���e��m�r��g��w�GGsn�������3��G���@c��ϕ�3k���w��A��i=]p���#�����\)��K���ؼ�SC�w������X��+9�����}�'�az�ƛr�+%"�|�'�'�c�0%Bk��6m��	��
1��*��_������G`ز� ������D12v�CMj��o2�������D�>�0 2Px��U�f��Wپ')U��=���@ՆO�F��>F\G��" �vq^��d�Z+��;<�F�ږN��lq<�����U�
����S����S���=�$��3Щ��4�����/g���p�\�w/��d^?X?�#b��*�C����,�L ��o�>�՞6�c��m,�������q�����W�"lJc���C���Oĵf[�|�@�G3�ʴ�]e'L��ʻ��bH��t}�Drl]���"=UV{�ʐ|kW�?�Ӭ��I��f���cI'n.�kC��6�J����˙��lS����������g�&��1���������$��Y�S���2��i�a�&��E�4�fz��������i].�	Fb�d�/+2�iO����L��:��o��"B��^C�	@�ŭ`&��j�ə�v,���'Ǣ���xL3	i�~�������uWY�x�)P~p㭳]&?a� �8e4?�1VW�]߱a[M��d2��T��fW��"95�k�_�^��H*���SCG����|Bcz3o�������O-r� M�F�C�?�?\�li8^T��~v�:�u�n�,�
�R5�o�V��ʙ�h�'q�N���
�O��⋊�z������hD
��a�p1R�"
.�����>hP��>Yi��y��Z1d�W`�ꎘ��@�N�$�����.'��Z����M�db�Y��t��Ah��7���T����s�h!����=ef��6m ����F�L	��9�0_ZL�@~�TbU��\���0��n�hB���8��D��h%��H7,��g��fE�J���?!����t{̛���[*��p�*�3a���B;Eh�L�'ø\�G��.�$�f� T$4u�+�5��}�<�Ӛ/�^��v* pBPS�Ԥ7P��kc6[�x�;��k�	r"��Z�3�8�U��Z��Bꡒ�V��dʹl�w��'��Wz/�zh��(͢pl栆���C$)+0����c���f�R�h8G�TI�Y��M,��X��|20��XN�nV7��Ľ�M�F�rc������ �0R!���ܛ�ݧ#6an���L�ɱSg$�}/[���Yv̄n?�T����'T���e2�s�0�@�rq�>;[��3�O_ �\P�Psgǖ��?����_�<����1MAPޛ裤]����}߃�Ah����,�O`[3.q�MS�r)��8������l�+��:�L����y�!��� �+��������ӫ�7=O���Aq���0��f�L�^Q�>6���f$�oυג(����~Yi)#���;a*�Y���JA�ί�ȸB�{��sQj���p$��1H_���΍�,,����q��P{}-����2�tZ����G�b2ѩz:�b4$�|��+��3k��8���E�A�C��m;��>\'ؠ��t�DFs:�y�m���j���%�jb�>�5��^{b��A<�D=��8�_!�	��/��T�����JE�%1}�;�q� �����7�Yg�M�~Y����2H���wf�l������{��w���A���h����\M��+T�-�f�ct�6`z���H>|F�x�j|[����,��=�1i���>��#��ߚ��"3�����w���%��?\��;,7�$�=}4��_��K�/̑J�8=�%�[� �2���N��ou�^!b'c�B3 �l�6\�ϭ�&;�I�{�����1$#����,�[&Xc�1s���AZ�D�G���-��e�*���~�=�$2kb�5\�BiBη�ѐf!`RMkH��ѓ��V�HCL5YQ��0ߚ4X`��q�=i|��<5Y�	/r��,{|m��~�񭺃�=֨N" ��}��>n���k�m ��S�K'̗�R=.�~��z�<yw��\��P���l�}�%�tщ�`_Q���
v��o�XMU�������m��N*=w{H�'�����a4oB!ހ��y�z�_��?�,�#}���C�WTykN&����<u���d�Z�ͅ2tB�!]_s�i�A�1|��g�`��ח�e��@�$��?���RW��M!�π�e[
˩b�]IVsa�<"@>�oО�� F�HeN���ݲ��P�8;�x�D�큋!~/E0���޳J'=���/��p��Y�j����0��]���#qX�C��ԅ�N(�tv!�s5�\,�<����?��B̖>An�B۔�~�
�j-)	�s�C�9/Hhv�Ɗ����h�ܿ�Cx�F�)UG��c��6���t�?�͛/+��6`9ۏ��e��4���1�b���K��/��?������?�Y1� �Z~y��8HP ��N׀.B�:����S��A�z@��''��-N��G�:-��c�$���4=#���D��NK��ҿ:�"g�qA�qw�+�KqB�`��Q�}Ǭ�Nۮ�i���'[/�dFe=� Bv ��ƙ��χB:a�[����𴔾��@�&1�D���b:�n�uTS�Y9�v��!�+�f���}�Ų �$,���9�W�L�˷��K�|�����O ǇG6����r�%��C�@�ż2��	����E�c�Y��]{��T��瀁��3<>�l����{) 5H]֐��ZoK����x�8`�f~��>{���Why'�^����*� +�B����x�qi�����e[Z���ETO)5T2Ys@H��7�)��wv^q51�@=(k5�
H�{�;r��.E�JdO񶸻6�bB�ii���������A�{�I��6Mv���t���>�U V�i�X8xćހ5^�A妠�-�2�r��v�6�- N�`Y+�k��!���nȁ�_zwm����aVZc@T���ڥ��鵿��3��|��hW^�	��2vtM��D OM�Uޣq�&de�n@�$��rVc�ڢ9]՚S�#A;�5���ͯ-�w7,�)��w���=wpB/mf���G�Κ��+7�xE8�a��&�0S���l#�H�2w>uaW�������ȯ�H�&	J=�@%�	�$,�?�Y�9�rl"W���o�Z|XƿBA��]����#�=��x��*0x��6�-�J��?��=�T�A�X��P�y��:�[�ȼM7����hp=j�%GH�wрK�{�uV�d�����	:Q)��P��A�� ��6��B�����e��4`p�Q��'s*�zB?��4��ܚl����]}�%:�!B�U,{a�g}]3�2*% �m�"ԲC���,7�^�5,ı B�YSYI��_�[_�h�13�I���$�~�)P��+�C����_U�c���i�%"�,ܽ�t��Ȧ��i����F�-�. L,�9^��2��#LY��ۻ�o)���k�@yr�S��'�='?S�pexd^���A7����؄�d�&x��nILl�;�<sX�7��P$�6K�ډP����t�2r�M�QM�:GRs�3��i���{zr�t8�-�y�3�S
���f%DT���O�꿧m9��$��n}\�#[*c1������2гg��r�7��t��ZC*�*'��!<d���<�A�9�)N�U�1O��{��2�:��<������S�R{��CZݹK!od����Y� ���S&�J�g��P�� ���f�~���1�B�Y윑ȊX*K3�}W�'e�>�r�VWΩlK���&׃6�B��}(S̨��aj�O^m������(qfc/#��
��e�5D�>� 92�k�֩0WY��D��u��6cɼ+�Y3��H=詋����يϼL>�W��O����p{&��m���q�����|N0V��\!2�JȜ�kAS-#x���!#gӺ��<~P����wmܙ:���:[�9�%��ʏ�A0 iMՖ*%e�i�>��<K�(Ap��
�����2��	�"Z�w�:��w�dC(�<N.���߹V��x!Z���W�|<@��x"���<a!��'��+����.�m��Hݦ�m(F9S��Zގ�p1S��;'�㷏����4��$|p���ٱ��{@%^��
E��H�Ð�~e0�����]��o���]�?�4�f���^�R����{$N�8�0o�8�k!���2| cO�}��$�8o�|��f�r �3����ݲ��$� ӟ�uoV_�s�3�!RG�;X���z5>K���Ĵ	��*�s<$�L ��'b>��;��x���e�0r#�@�G��T[?��AI7�g}���ԥ-��(גd�κ�>+Q\�>V=�U�#m�UVh�+q��8�?P!C���_��:���ͷU��=��[}.{�[>=~�r�6�W�LH���9E�o��y���2��5����k��������|Vk���D��kI�q��X�H�_:�MS��P�F��3��4y�@�K��"����"p���_�yU+����Ga@{C)#~ݱ�#�0lN%��Ke����C����� �y���%V�[�Ԟ��X�6SYg�y�&|՛%WҰ_�g�C��_���U��,��Uلh#P>>�W�";�F�=�
�bݎ���px�틵^�{zs�"RD\��L������}ըM�3|Yn$��9�^#^`������<���\o@���msI�����UlC����~7X֮���W�_>^�kƽyF��a�HNNb�UP������C����G�
*��c$�+��E|��,g_]j�<&�L�&�l��o�&��s]��0;�$_��h��X��<Kq��ǟk�lEZ�囱�h:�#�v?�X�mRag��CS5g�.���ĥ�{�9�8�ܲS�:,z�4��t�v
i�VC9�����,�N�5�Yx�a���l��Rڪ��VZ.����aR�=�W��a�\瞭D`���&à$ک=/ŸC�v������4}h��/H�m6{�j�D125<IŭVs~�O腍�m�{fH�a�,>q,��Q�wD ǵ"#�Q�EW�$uk����)�^9��&� zY�*����7���l�Ew�f: �pl��ϋrǨA�a�lk�����@;aD�D�0�!�q���z�?G*��x]�KQ�D0�P�i}��" �����\�"� A���5	�t�u����PHGE�����@�/���v� �v�v9F>��҇������@h�|\���z�bbՙ&��QRޏ갤@��L2��R�^�yow��Vq��M
�C�}�y0V�1N|�!�8^a��:���Ϳ�ܶ9[� ���ڜ����{pdf |���Rg :xq���'a��S+O��q'��[k���\���9V1"K�ؿ��λY�6�`��L,�N��Lb818�!�e$���/�"o7AT֧1�� �n�>Y[x��J޵����t�f8��Kt�I6[����_|6��fx�~Mm���T#+u�R*��r>�_�"ɗ�Phb�.�Ym����ԕ��@|f��ʄ׉s8��]֓�&��\�R�M^hy����,}z'�I�H�m�`��v����5%�7^���֏V�֔F��O��#-�I�|B;�tz9�ܣ�I9Q��tф���?n ��-���:EL�2�`2o6/��?X����&k� &�����מ=a�dM�ru[�q �`�R��7׉�	)c"o�`�9x
܌��=A�4��2 �'�~
A;s�O%��ߓ����rh��Ӡ\�9��<���~�cwY{t˂-p�>��ݲ����;��M�%ܗ~����݋��
$�P(���o�W�U��AH�kS���-�q�6�j��@��Z��p��^
c&r����nU�
�\�k���W������r�����8��db��f���r
�M�2��ѵ�,ڞ��1i����:�~!�L�.4m��,����@��`PB5��}���F�HZq�۸)����Pt 
�T�W��}����IHB�Җe��`����-R�{��� �|���v�N�( �6vΣ-��v;��4D|�����ެάl`�襲�B�?!�����N��Ѯk�q\�ڷ���H�\�*�&������T95	]�;�|Ǔ��͉=4&��f��"���Ӑ�hB98�n�����4�u�P�n�jU�7�����9l};f�ϑU��kFBy3L���l���7�R^ƔT�ī8��F'���ݣy�c,��]#�|��\D��A��T���F�T�Wf�P7��}Z��'�5�<�L�#@����+�$l8��b=!��
|�����5?�k�@��T6��Qk������%�#z�IL�֤�����Pw#�iyq� ZU�?Ǽ����2�O�]6��X���b�[읗D��q�Z 5���d(Ppp\Y��Z����R���hf��!�x�<�;�ǖ�9GE�(X��C|��ĕ�͈E�Ȩ���n��1��l�h�O�-��[aL�4�r|�g��MX�@YlϽF�ǂ*�]�&�~8Z鹃����6��+�נ���us��	^!����ə���`c�s
���l�Od۳��� +��ҁ�A�[�@��>�Q�v�9;��`�҇K�ʣ�_���¿�v�����!+\�O	�9�RL�Bc�AR����'���������%觏xT${5�y�ycQ�v����k���BBm*ئ�=1�u��̀�	(�Eil��R��H��&��3�x�S����>�Uv�ބ��,����%�s@L�)�^�-��S���ӿU�=�1�	���8vǂr�l�hS�>>� x�T#��H�v>�独�X��B�Ut���]�}5����4ixz~D�n��)5˘�3Ȇ�oK̳�`�1	ꉊ�ɛ'�ώ7����-�l��ɬ,LtQ��E���pSs�;���-�Z�0F�)n�&>�=	�ٿgn�^��z�#�_��n����$��&���ߪt���	�����i�������w��T-s��c[6�/�t���}X�*�۫���2���"���p��H���e%Q�����x{���PZ �:��c@�����ʟ9�h�O|[pҔ��0�ӫ�Ќ9Mg/�./�h��������M	el���#��'��?G�,��ܧ�Ŋ�~���4��4������#�^5 4���i��fK�N���ɖ�1�w�����u+�c�g쉲��Eg�:!�16��Hhg,;F,������'��}��,ijaZ�<,�|e�SEN�Sn����Y[a	�ay��	X,��� ��� <��C}�#7����2#������b��OA�;V^�N�U���z]Kq3˸�&�U�M	[W�fU�,�C!�T,;6�")�-9bC�fj~����-��j������brާ`"��2g���V��vj6L6~����<By�G��R'?��������m��5�_(ݐʝ�iZ�܈������F"���#��gnq�?2�T5�U�sT��5��>˛�TѕP�깕��X�O���s�0� ƿ}s�O(=s��ؼ��o�V��NUH�Yk|���'���`Ar;�!^�K��=�э2�:H�`�2O&��tG���C�v��vU�O ��1��ͅ�F7>�}���z��E��u+��,�]��ʘ*_�-��,#Sxˍ�ـé�3s>P��o���Qm��$�gef��#��Q�J�N�����K�lg<�h��V 7�`Kȧ{0"?�˫���.Fm�k>�	%�惶�g|q���{~6s�Z��nM(S�	g&�Oo�&٥W:��ꋓ�����x�_��tױҌ
�QL9�n������̤6��M�S}�{ЪXh��2_�
�'��F�b(�Js�7�Jr Ͳ�FХp�#:��C	L�'9�g��N��˫��>R��3�����\�b�u�Ǘ
H�QbZr݃���'4��}����� k�=��A4m�����Q� ��G���6/��J�Ptĵgn�h���m��[�¼�PD���J ��>r?Ut���۽B������!P���u�q(��4����%NQ߽�1A�����K�;&�&��wq/tM�^@�(O�yk� ���r��Q�q/Gw�����XpQמ�U�U���m0��BU;�
����qg�����/(�5��u����8�a��y?(��^�7�u��d�Y�|\��Ţ��g�̠i�ʔ6T�}�b�jGO7��1��^��L˂�����p_�͎��V�5�=o)�N��|v};��0!���H ��t��W��Y�l�3k �L����މ;��3�Ŏd����F���6�@�"#���J��ʨ4Y��)ݳ���\^���ѩ��)��5H#�_�x�7�pM�#�4��O����L��B���y���#���5�|!7�%5��`s��R�TS��=�Ѷ��8{̾A#?7.��3�z��b����x�灴q��u݆S���!�'�4Sd����X�.c�^)��4/&�
�W.U�����曊"��YДI����Zq�)2<���hLJz4�$�,G�>� �y�ϗ�� ������^O��>PB�ԟ�]p�6�ߟD��Ӫ�-`�V���;,��}��y$J�I�QAÖ�~[���n~n���գ��!�ҍ2�[F��gɿ��v::����_E��B*F:
��#s��U;C���Jdk��~~���4!L)��ҰW�$��0\z^Z�(F�<)�Q;D�V&�?��>p�R�8�Y/p'I$B�t�	�>����6��og�K;l���}%�I��4n��Ÿ#�A��+��Fr2�^]+�8�7~Q`zш���M��m`Mec̆�����ja� ��O<��~�"n�8;+�5�0�n���pcٰv�ױ�s�KCvf�H/I���@��I�izʴ'Ro4����a��&<�(<1eL�z<�����e6|�<����)0v��$ ���
�Wr(�V��sH�� 8EWsM�X6�:Kha�mf��gG��I�V&��E2��@Ēx�N�GH�#��DX������!����`/�����!�9�'�rY�$��� Rc�^Q�.a��;I0˟����y�[��l�������P�P²A�l�����x�:�':iY�yo0hz<����?���'�_t�9� �P�����=H/_8�aեo�d��DS��6�F4�/��_�s)<'���L�)E�qD��3?��6�V��ET�~m�__�w1���̔)(�
�dJ���G����<�"l�4ٹ�G�T�J�����V���~,-�Q�x����E�4մ��n���Tɺ�7�����`�3S�fh�9�������"���@#885nOJE��p��r/����u��P��R�.Hc� �L����ڥ9��}��Y�Ϭ<��v'�)���ef���7����jf7����>�!�Mu�uDwH�^�1��A�+�3c�Lj�Hh0hw'/�A�q���ɗvk��+Vb?@�����*V��P�ѫ�,U�VD�f'w��c	t��JuG9M�AO��]@z����6�ʹ^����t��O�s��s��w.ٕT�^��?$7t�?r� yl�:O$}�p� ������US&Ͻ�^@����'�Ԋ	�~��I�&�	��_�+�ڗٍ"�<�5a�&~ϟ��\�����֫y�w���h���vZ�-�\P�mm҇�j�*�
 E��|�`���C3�z�YY�7����S���3*�l'�,v�L\:���L��vԁ'k]%Ӌ5�~�
��He�{�3�khj�A�A���#�FI}�T����fvDC��׳�*�_��x���6��}_���m��"�s��uJ�{o�����@[ԁ�	�3irJ�yқk��J����m\-9]ś��� E�Ǡ��!���UIHE�Bl��%���<]�t��~�9τj�\�r��?�%�ss�c��+�κ�����ׂ����8U}e�Z�kᨾ�_T�x$J��ޏ�ð�#�o9[�;�sS�L��#]�xH�5�#b��ԃt/s�gk�����Ȍ�l���2�m��_|������3�D\��������g��A�'�`�<���;���%�-ːq]ԝ�(�qoHu(>Y���2���s��F�b	��8�3p������ܣ���d�_�ȁ7֓�f4�ľ{yhH��ر�#����[�q�F�Tοyn������9�����v�*���3�7I:�&�c�5;�|��v�����0 &*���_j�{���"�h��&W�E�3I2WrX�mj,��-m@Q�����e�e(��	)��:�����S���֣W��}��X �FiG���uӡbt���w�O������ɤ7�� j�{u��d�|3vC���S�S��H�T���[KVS��c9�������h*�i����K���%��}�Gڈ�;~/�� ��:�4l�2���3��^�YͥW�W�x���{�Tu�;"|z�6��$�SWx^<��+NiQC�����q���������W/��Ӄ%�z��;ݯ����D8�Rγ�pTwɣ��)��`�I�F�J�"-�����ٙWE\�Mk��ކ�������5 [�ѹ*����1�qă���o���O���-�Ph�)Z��SksUQt�;��.{k��}�FZ�i~�;9Ùݰrٟ\��:�kg��� �>-z1�� 6�e뀄����*t��y� F��W,�B���:��Z��ΨwY[B����
�Ծ�lʷΦm�#��F?����C�S~M�|8O���,"lʯ)��y핆��Z�T����ݺ}>h`U��>l$��9��4C�4��	}`{kE�<�g��#	�w�|6c�8C��ll�n�s����đ8?GbL��L����:'��{
��� ���*�z�Hs��CaÏw����3}ij�P���A �%|���Pxݟ�8I����_�%�KE�T��� ���7�k��.B�mt�>�XPe^��Jص'��#쮏]3�@O3T)yTٕN���6631�F�2U7s�9� ���~Oz��d��"�C���-3�u�a����g�)Fj�!N�(j��1��R2��T�ғ��F۩�;��؍�UD��x�E_�m0�ބ�N�Di[��N�X�xh������;j~\K�>
��.��>���'Tq����h�E��>7����a�PC3r�s2�'II����V5��X|}���@9.���A�F����ZHb��kp&G��P�B����&�w��\�h��*���V�������,(�Ud� zZ<o�=5&������̾�j�hy]��c}�h?� ��7�iE-�a7U�׻i#o{�v��)b����T�Z`}������/�i�^���L�E���v� C&w�S���ϋI~��;�o��<V"�bf�OZ��Ûi���G}����$�/p�fڷ��~iF�������e}�������[K����v��[��E^���4�H�d�|�		oT� nm%};���jPAZv�!�+��m=������:�~g�2��Snĩ�9�,J. �i�j	��i85�V:��%@E(��}�kro+H�����L/З)��0U�a�&{@�`3<��z�T��Q�1���G��'�R�@(#��^&��������O��i�7C�����OHj�#�t����@�A��'�T\���$�֒ȣ�q�$8k�5;��2&F���%FP\oW�p�@�_�B�{ɴ�6 �U�gQh�]�R(�����Oy�������@c�3[�M,#�>���{�%�wK�I�.�v��63�)��.&���;���?��g���5Ζ���S��|�w�A�m�1�^�$f�f�Ĳ��d��U~׾n*Wde�[a9��Ĝ󱞷��22GN�|�qsވ�p�C�VRm��A�u���J=wZc�u�[Ɔ'C�-��h��:'�ڒ"�����!%_%x�=��wp�b
(ĸ��=e��ȏĲryIp�ߦ��8~x��Ey�c��g���@���ݦ	�9EgұN�\�f���j���@5�e|�L�V�H4/5�gH}��i���D
���~ۭ4�=t��r�� ;�!��8[֡����e�����7z�<���߱}6��)���zd���Mߟ��YP��S&��+��m�8�̀��G�}�rQu�Ј�/���i�pp�����]^��]��ǭ�^�ښ<�%B��`�ޟ�s��M(-߾܂�[�Z�z[x�iG�q����i���0MyC��d�
P&^cKy���@Hl� uf�Ӑ��"��#y�c��@����rjS������ ?o�x:�J
z��\�5��y�.<�F�B�}<j�R��n�X��T���§���p>ix��Xu"I��8Y,D%�'Ϣ 
|�Ɂ�B���\�����}�!Ÿg4fX��G�ל�O�+��g�O��B�@�g�5�VBS�	;��Ι]��!W��]�_�N�����$����ߟi۴�iE�pp����q �)�c�yk�H�ueV7̒p���\��i�g��Q��}�k��Eu�~B���??���@!ְ��'+�2�ެ���~(�)�X��+%^�Fy�>nlLj	4�E���"Dp��_�PC���f�4�ڷY6���g�i7�X��[�]�iu���>*�Hخ4�����\���{�0#�^�u.�r/S����������G����׻��ޑjebbx�#����:gi�ǩO��Ƽ�P�9c
�p��o�Gk�������E��&��?�.�N}8i07R�$+>���\ꓼ���6fy�$��e�@�ܺ(dK��yy���[ٟ�Dxx�c��@����ֿ���S���N�z{/����rU\i^���!"�u�����/�~$���*y?��h%�����\����}[rL��;��63� 0@���I>Op�m+͎��d6��T���g�ʋ�Z��<���"L��'�'L�| �pS�51i^a��Y]E��&pA�.c-���mi؃U����?;9�ߘ7��<a⨨��}Yvu|�l����|��e�]r�%��5w'�]n��9�\g�4��|⪝q� �L��ܶ���ÒҶ�[m�f��Ż������8+m=�DJB���ҿg��vv&���4a�½�NU�i�D\�1��G.Žl>|Y������>[ŀ����������͌\�O\GVl� �}U�4���=��Q�z��v�nC��5�\͐jp�{ ,�Ҡ�Dr6��s���]��"��$D�R�����G⠩p��b[G�Z��M(>�o/Xn��25���9�e2������a��n�+E�pk(�)��W�%O��i�	!���+�oܷq�ﵞ;xI.����6�c��)�:vIJ����|�D��9��HP���uC*�O�pR��(9&�G��]�[+�xZ��i$"v�z��4�Ǔְ}�sW����T�y�|����a8+����@�h�[���E�GBGf��{.�\����Tj�Y��WLjqD*R�u;U	��{QFV�� s����4�����ٻ_ʹ�}UI�M��.3V���eGѦ�F�V)����$V�R|gq��Ӎà]���5I}C&�_�:K]`��^�����NJ���ŷ�h�4Y$&�W� }O���K��Rg�f�{0�tn�&��u�D(R,)p�^ޙ���99�^��o��m/��gmސ�h���3+�B���{��v��Q�����Q��d0�}0@���䀯�\�.����_B�2�^K�ΊT����Te�]s��,�:D�zM�L��u�ͣ�
_ T����e�3���0�������	k���� ����L|���V���	�[a9�w���r��O�A��{T0��Z�B��#�d�&7z�1��B
�X��lc d���q\F�SJ�_��ǘE�׻�R���>��k�-����8��/�$e*�p����W�ofɳb�S�ɍ��bW�$�ǫ�z;$V� ��p��hX0)��YVY��m9I�^6�zzQ3�l4;���e��Ok��-���"�#�SaE(���Qs̶�Y�z��J)N3�K¥��#e8pǥ���߹�}v��v��"@-���;�|�p�>��Y���C��j߇�U=#�{��<�^�;ZaUy���)�@�O��WL2X�e�a�szx��I�7ֳR�_e���t;k��Y,(���8�}��Yxfo���*���|Z����Qrs��:�O�uݪ��d�XBK(�fv��jb���,&���[��5�c�Zյ������f5�,��c���x]1���~o�-0�Ǒ�� t�,n&���b�U�Y�Z9�<Dܔ�zX<g��������
�0c`$�{^��?0Mp#�=��}�l㙁$u�UC��an��������	��c&o�4��csy�.o �Cle��ZQ��9o)fO�`+zo�����~�R���rZ���x�sw���iHP�'��?��-~�U��ڳx{���OT��Q?[�}�y\���8�;�Vc���nP��'M�s���9����!y� �9����c3<��n%�2M�||��|��� ���@�Ǥs6�|�o���nV���T��`;S��?�VJ����".���)�E�!{��uڶ)Gaq�o�E3��1KƧJ!@��ՙ�
���r9������R:�������"L��&����
�uw}_��}P�<�x��3O�P���`X֘@������	��$t��kq}8֜#൒��Ȣ!'- �P�D��<fw��7�&�*��蟔�U� 73��|�Z��d�?A����U�����,j
_�\�Ǽ%����q��:�R��}9��g"�'�`�3+xi�(�Ӄ��"��ЗB�ѪI��/��\?*�;�J�w�JDȲ6�;�*��ݕT���#������&�K��.�{�)Nsaiè��4�"w���(ġ@Τ�����Z��+�S�� Wv��;��̿	)��g�Z�>N��]N|+c&�!;	4:�����f�����6��6���2�z�����}��))@O4�l�3D$�T�Ѽ�1��1W��M�c��"C=W�V�7����"�_(D�j��̇|���f�yn|h�����ط��ő!bI2��ؙ09���,������.��Ry���6�-o�U<ǐAo<Al���(�'t7��@�[ت��B��~v϶E���,�3�;=�ÌV����z.D��ƻ0wC�<IlQn(~b;��g��)
�r��~�no�|���S�o17��pOY�l~��w���w��C9��¬=*��Dr�������{�s}V�[Y���6��S�m�^ѭ�h�q��ٍU�����L��Ddڶ��³Z�i�#zOF�b0�]�.j�+�I���F5�}0��y.y��� ~+�O�,KWD���[�5��|N7斎����P����+&�
�����6<K`D�v��MKϿC��Z���Y� "��	�Wzb�ѡ�0�<߆�8y�4a����t��J��x�$�
E����B�M��R�!�7��I�����K؂a�s*9�n��i|$$go���Լ���']��Q��ߧ~�*�����J��r_�I� 4'֡�Q�9Ԣ�)���7�.�3�����*���'��\���9����,��#����Nq=����6��kw�7����̈́$A<�l�>	�F�x��+3�����F�4�&��Q��M���}b ���[�s�A>��Nd�'�s$���?S!������!d���e�-2�F(7��Z|2RT+z
m� n�ċk.��a
��t�G�eٞR!g�����U6�f"��7�}¤�iv�uu�#?��)��s`.))1
?�Y�j�����xܮl,���K'�+�uz])��
?�'�>1:�IS��,�o�;�=�sDx�7���c�#y�&�"�!��>�=9!0����K�~[5CŜ�z�?b}>�[�A�'?�>� D�J�sH��q��&�c��]E�	����_���N�>�ɒF"�����1R�w��������۳��@�p�����Ay�$k!���i6�3OqG�!�.j_d���-��{Gp����-���$�n#��[��C<��4�r���k�p�Ո1,�yw��*�Kۥl1N	.�\�b#�}oI+ �7_Sv���j=�P=N����rw괡���Ç��<�jP򹬴�I���OJ�g���J�ӆ:�Z�_+�����:86 �Z�90p�Ռ�8@ԇ��_�]�w}��R�v�.L[���x������u��IQ+(�7��N ���'H�P��~p8In"���`�7vא�7���*�H�q�5]y�g�pv��s%�mA/��^K10*��\�Ȝ�#�O�7:�Z�/Cc��"���\g�b��]6�"E�e�� �&;B�>�H�x���$\�$��c��S_*X��P\@Za��sfm!�V�x�7����
�[�w6�8Ї�͏�%���f��]��p� �6����閬"�A��u(p����!x��:-�U�ˬ*| �}����ʓ��&g���a�_�A�4f���]�����4���ɨ�?�rN�0�@X-���¯�1`'²��и�PC�O�rFD"8�wh����k+�1��$����r�!jF���:��|\j7Dse88lV���]�QB%��y�`d��p��)/{�V�y � ��?���Bͣ�xS����h�P[s���Q��y�*�w�2�
"�¾md�1��̙:�(zԷmO~��by�W���g�B0{��w��?k5�C����_S�:ğ�*��40톰ʏ�P�!H�\2x�@GT���^����Q*¤2��{���#3�۲>���=�'��C�q-X-g�J�X|r,w��5b�k�͌y8Sbx 1&��H.�Oq���?�H!ؾ��a6?����j�p��.|׮-NѸ鈄�H�/"x��%�U��ʆ�V-�7K���FV{j2"���f��ī��]��F��o��D�"%	�#r	�13q���a��I {B��.%��|����)�\̈o���q\��+x K��Fu㠓��Q���u�煀�����1�W�1|�˼՛s�<�3�>�CO=hXJ|m�zW�)s��ɮ����:$�`�����>B4���@K����w�L�?7-2�+0.��U?8e�\�Xs���d��� ?���$����N������%��VC���N�G�9�;m� ˒�jk(OP_!�N���z��m3�s?�e�	�<�i�R�� �@�ӴǳA��>����(�dE�.���1a6�/��w���Q���(�;�I[MfN�M�V���%��xի1×�o@D�lkU�����3���NW��K�z��n]cm���;��΁<!�4Җ������B�D*'y�⼹\g�_�uz	�m���XI������c1GpQ$��u�c������q�4H�mހb���J6���7(�Ȗ���i�l�� ׽����=��xų�OLD�v�pp�z�>�J]�̏#gҕ����cu�����3C���a�6H����<�6-[����' 	���;%|���YF��wK�V�ht�ej�r��@��1keJF.h�.�@Co��������H�v�
��V�m��P���m!��2W�b�G������	��g���c���oZ�#Z�椙};N\�Gt8�sI_��G2%��w��C�M$nI�^]2�-YO��B{��^��!\��i2~X�_��>��Y`�K2�2���%�+ǁ�R���>8B.C7�ȯk�����y��G���@5��������Rd����>Z�� �O���C���K	L�~D���Й���5�3��X���j�m���>Yz���G��P�_�1���~f��|.-Q�=�*ZB���L>�����"�@=�H�\RQ%؟^A�����4e�D�Cs��C(m�����!^�.d��;���	���'YerF��sua���PZ@�4)�o|�
#��Nx�Op�ڿ��y�ZK�𹤿~��Ghz�&�;�0�����0�������Z_jcX��ͪ�;��6OJ����f2oC�ϰqf�a��b���/>� &b�12����D�MH:�X�������#q��)�V���}U�Yd���"W�> Y��I�FC�G�2z]\W�7;���}4�Z&���Y�h(��AO�܇<�u�*m�C.�\�az���
��d-*Ns��˓M0v���5T�Vzج2٭^R�)����l����7� @������iT�o�����JAF<���^�j_7����ꁻ�0������C7!��
[t�T���}H4	L���~B$�Jrb	��ĉ~\��J1oK;�6��{���0)3�_+ⴃ��\/@�G�'PxY��W����Rj	"�^�1C]�FD��]��V5ҹ�����*Ԭl`[���}��:Ux��h�v^���/rm�	X�I܀�t?�o66cq�˷ds*�����bö��p�K
:Gh�bޞhG��W�������^�}��Q�"B�����,���n6����`F��;?c{޺�Ū��r�L�Z����åW_1m�u�y���i�� 4�@* w0��A��H��0��6Hb"@|VG�K�c�����nleyH0����;�2���s#��إ8���4���5Q�悅{��W靉/8��w��&�8S`R�>�g�j�c����x�ɾN'���0�����E��o8�N}�Ǣ{��R'K�Pv���h��P�/b�ݎ��c���F�;�J���V4<��'�7�[�+�yt�y�>�Soi'�`_����u*��&c�b���[Y���{�����p��bQhB-����\�g	:�Y�3�w�eCSĽ�"�Q�<$)���b<7m����`Fs<T;�l��(�L8��+�����HmVN3��R`�sqB���N��%m ��nŞ5AA���2!9_3��K�F�_�#*T���l[Kn�,�����cH���4#rA.j\�FeJ\�\�a)�p��U�3JknSXɜ�WD���6�M���W���NX޴#�]r
�-�{L�I�����x��ʑ0Ӿ��Q��8"��%7��k��&C�l��E򏮧4��]�UA�k��ċ/CC�Ow�`�4ɚQ�=�h��L9k\��bk"�:jN�����QTW�P�F���4��Y��:&f���M-ͅ�j2	�=��ZH4j���W!t�,�N^�Q������r.�O���ʫ`����Xt"f�%�L�}W�a_U5�Ya�{c�6���q�"�[�c��{m�N>?�~�z_��D�D����i�si���.�b����Ơ�H�XT��H$`$Y�l� ����|=V9OG2��4�ʏ�~�R:N-�챢=!��f�	U����^e��d�Z�ty�!<��־ai(?�cw���F���}�hc��b��,d�\���N����~l&e}��ɺ]3�W�䃜u�C��o���=2$v��E������l�K�-����aii&W�7�w��L�X �,�����P�����)m��oZ!�g^��-�H[�N��\a�s��LCL�
����H�n}����N�Qr���À%{M6�����vqI�V'ԡ?�6>���k������U��(^�阪�3z������׃b�>�/=|�Vj�����L0A�F�G����W>����f����{+�+ŧ㰛(����(�M��U��%is���MM�����Y�7�C�� 	]Ȳiq�}��jgD'�C����U������<���������Xp�E����5�xG*�s��ĭ���ԁ�kZO lZ��'�[�x浆ҧb�L���ϒ@����_���hw��7������%�nb.��(��eC�b���|EJ�2gC�8�Ss3��%�w��яD�%=�p$wk���D��<"�?2'���'A<?'B���6���F4i9�	�l�8w+=׈f;�ۺ�@.�S��㤼�G�1Pjq1����Yy�
�)4��y�'>��\ƻ�W�\��~g��r^���������^o_ߤ��O��Г���(�	5K1i2]��q�
8�4�x��Dr:�,]�i�-7X��[�z6S9����{־52�H��f'�����V ӣ4Ӂ#�be؝&)��Y[oS.��=�#��o�Z��X+�f���e�S��ℐr�o���p��Gmf�E��]���ɾ�a�c�M?F����� ���h���٪ �#�{x���/���<������<�L�$I��
�p���$���,�\hF5i�f�!TU!o�7Y�d-�:���Yy��-)&���Q�&�d��&ev�;�'p�n�1nǘ��ڄ��R�B��H�F�~���El�r�`5�m@	_���(���Z���2(��g�	~Aw���
�v���+w�{:wg����~-�hYV�������O"Q�e9�~�^B>30��0\ы����H��8�hR���Bʭ�n��0�x!�k9�I_M�C�~����Ѹ���7�ݹ�v���=!�o�8�~}�S9$�=Z̈��5�ᄌ<��m�n�ps{�	�9ID��<�'ua���we*P�khO8���1�)������7ػq�2�}���F���5��~7wcC�9�Gi��=s�j=]H���E��d)f�R%�s*l�������?U����vo� �!-��"����D)'�����frA����k��P�\�3�k4� ��O�aL��9$�ʻ�.�Qb�1��<%7�O'�>k�2�ݩF�;LD��'k�s��1+��C�0y%��w�o ���<��y�����³&��D��S��s���f9x����z-)U���[���O����Q�eb:t�3#g�m�c]��d�� �{�[���Qo:Zi%��/�Bg2�ô-��߭
*�L�=�������kF
��c�܆*V�����9�z���&�H���f��N��+/*���Hfx1]�����ͯ�������@B>����-���X?~������d���F�&
U?����p��q�)�M����+R��29�FH[�|�.lq1Ap�^��X¨�Q�w����챀w��U���U\��������m��0��i���x,U�]���:5�+F�!��¥�|,����~����=���t�8�i�i���~�d��H��]��� �Q���ѳ1R]��s�T�$�2��ۍ缇�'�`�*������k��>���T�b]��W�At�x銡4>�28	��u""�M!%��3�õ�(@�O�7�M�L���|`��b�7m�����������}~	�����4�j;��1휚Rl�,�EzG�)��FLy6�>����G�6i�4�����{Rf���Dl�W߬�����+%�%����h��9i~��[O���-��}�X����l:,\�&�*fp�>Ԡ����8ӂ���ev��&[2��W&�?Z�"l��-�qFx� �Y�ڽ�^܎d�a�Mg!c>��.�s^�Ol�S2,#����w����8R��L�h����3�E��.hNr-���)7�G���VB����+���g�G��w:KI�����^J7���¥�NWv�El�n]�4��g��9&�����r����x`k(>���
�������������\����Ͻ2���������L�������6��ڻ�n	�u�ݘ�u�=����Nw2�r�����cNW�����gzo�V���,�.M��?��52�{۾{K�_��o�pZ'��OO;T��� ݠ=Q��j|�ͷ�ch6F@���H���se��t ɇ��h^�����ܫ�8_w�N�~%��-v�Qe����p�&��Ǹ�½T����f�0�Ɏune�P��B�6��%:k��I�����OKN.ǫ(��7����࿛xsF'�_�|�[ �+Ә�+��a����=2�q�w>��y�c@�R��a;k<m�w��x��9��Dۓ/�����h
�G)�f��	�%��0SS��9�1��}�����nW;XGi,ANZ�?����D^+�΄��V�Bm���alw��tH��(RL"ohʀ4�R����i�
�j<�������X�Z�t"uƺl���R��qW���d	�<�����]���4<���=�B0l��i�QH>�&:#c	:5�Z��q%�۱�K0V�}ץ�Fo(�$�lTl[�.[����	�$[g(���N�}��?�g���n牑&?�T�*P��No%���!�^/�3�����xt
���rsب��l��H��c���;�m��	]+�z�> J���(��_��	6��'�>�X�)����"u����~Cj�*frkۡ%6"���U�}ɒog�����?�r$!���m�DÆ�^/>�r9��mL_�<����
<y
I���n}��"������b���/Q��'$fk��"#f�G��v$mr�;�jbHņ�]�W��Nκ�B��&���K���v:U���0"
��!���̍�i
�[��%F�@"�2��;HU�1��K�yya�M������`ĵ����2�E�������'����q#�������	�r+7��,�Y:�v�d�go������^kr���eu�0��́���w��]J#������u� q 7)�]{ {p��0o�w���qI)�,��p��|��L��Eq������̅"���_�ѿ���R�@�!�+?T�*�~u�>��~h}j��)1 O<��?�D���Ѝ�J��椪nnQ!ќ�F�,$U!��6i=�ܒ�;��̉�9'-"��:�=���'I�͛��G��g|_N=�m���J;%�P������g�뒣>��{�G�#B���<
����aM)^0GQ=�婺}a�&7�����]��c��Bl���mOD���5�Uap!bWv;�Ҧ�f�����s�p\���|-�a	�I:���g�[q��j]Te�r�.�� dC�Z��:h�Bœh�� 9��K�NK�oL\ɢ���y�#�O!�Tp�������3���0�S	�F # ���l���˶I�����dl����`��$�N<+:+��L��fF�;�D�%)�B��.":�8��ђu^�v4:��n61��c�0⼁ٷ��X �ҭ�>i8��1��޼L�Ӄ�Gb�r��ʇo��e+˅?�O1�sy������$��(FƘ��öÀ���-&��,�[5l�H_h؛J-8	T#�w����3�����e>߈ña��u�~�o�=_U�Dm\@�~F6���=�w��[ w����n�~����T��՟�cKҨ`"7EV����6A(�:���c��m�q��i5&�J�r�����$��ℼ6����o�Q?�WTQ�g�(�l��@?P�jg%�a#�@���>��*[fy.��r�Wƥ�-#�A0_*�Ԗ^�s]��*�s7�D�!�cK���9�VV  &��*l�Q�����i_�+��4?۸D�%���xe� 8L�gs���߀":ڼ"��J(8&v��GƏT�b'%u���Ц0��v`o�NGh0�N�ٟ����lF\H�L����>����A���)&��
K�W��hQ���M���z-q��W29�Ն|����~��9�!."/M��qXFԗ�bg�ۍ>�$�H�F� R_��MC���(��(d^0�Ҥ���/�F�(ϻes��HʉJ�>��R��Ef�Y�����#Ѽpz�b��"��i��eT��~��K�tP�6c�k�Xw2��X�S��cQ<P��jF7t���io��GN�.�
�W���f���Qy�'`��h��]��!��`���kM\�;9���D#a��^���؎�|s\t�_��vԾk��ߢ��+d=�����Z�x;����ȷ��ٽ�_��%@�����w����=T�����Y�`:ow�u���k�хAg�������!U�T&T� �7\^�?��T�UQ�I�ʺ�_�8d�@4��:%G9 '1�T]����i�B�ޡ`m3Vz�gGK����S% kfk��l-I9�]��*����W���7���-|��Bw� Uk?�ɶ0�6�
�7�S7l� G���_���	<�Y�Ȗx;��-[d&������^.=����.���%E���c�y��i0*+~��D~��K@�*/RH�Z�a�2��h���VWO�\�������Q�Q?�vJ�C�2�`�!X�1��� ���ghК6 ݯT��w>w����b�	�o��ƠB�C	�S%@E��Se�cQB��NGW9n���P��x�#�M��\�ƕ�����\��&t��U��I��^��b �l�=�v/x�!���nh�e�d�%C�o(��#uM��Fa�s�H�?ڰ�,t����.4C�~X�/׫¬�맯xꁙ���n��x.*x��t�#)\u���by紏�������O,V�n���g(JJ���P{�"LᨖΦ��,�$.��h��\�9&qbA�6Rn�80�Ɩ]R}ڛ0�]L�#����Ϋ��{+�$A�A��B�\���.�ՒϘX޸m}��Z��(���� [m<}�J��:�����W4��|�Tl�A6"�}8��\�*޹���8'�N����t1��훞8_�[:\.�&��\b03�"����<�C�Yv�?�7�3_���k�;F���%��jN���`,�c_�F	�vL�Dm?	~`0�I`1���o�L�Nb3�1�7f�j�H�����@���Uc��OUnb�$t�XN���`_�+c�����sLُ��cZ�\Õ|G�L/�8��t�*VW���k��v�(��.�m�. ����.�.*��дy��w[�l�#�jO�v��[�o��T�6���H��ܾ:��`�m>�
|�R?Z��?z:LZ�,��q���[|:ٛU�F�uw]KհŔ�h��Z��w+Ϊ��^ei�ѷ�URf���}P��;�^f�Z�;:�)|e�l�Il|�Y� �H�H���]pu�}��պ���4���2�=au����|��IxgH(ș�<��b�Ԓ�k� �;���F��ac���?�e�0��w���Jԥw ���N�2��^ZR\\�V��YR�O�&�ܾ@��ǔM���ǎ��6�aA?7��Ճd��j����٭9 0�6��ͧ�A~R	� `�������'$;�jN,AzO.��X�׵Ͷ��'n�:�N�����Fмl�ͼ�