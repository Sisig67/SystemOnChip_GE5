��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%���J�(J����ؑ���s�G8*��\�t`���^2Jc>�a��M-���-l�lt���BH�`ߖ�����r=?�ܚ0B�!I��5��,_��z����ƕ[�hrs�� ���B�Da�k� �%�8.���7$��t�J��8�� �*L�(��L����D^Κ�'iZE�R�hSY�K�9���������v�:��K��-^$0��DP8J�@��W�(����]�NnZ\��R�)��i��hv��W֏���k1D�6+8q��s�U���CH���EΛ��~T�cSq�yثa�]ޣY�����c�Bۯ9Q�5���h=tI�E�v*
��szP�c+�?ή�^��䝿��8{�I�{є�`�T[�@P���&P��k�R�=R��܁�#�ʓ�+|��ih�I�&�i}�l�tjX��A��ä,�VJ���d���Ը3p����!����V�n�K���A�[n�sxe���!�y}�\�Е�X21K�L܆�
���0l��#]�k7i�j�;��i�-J	�v�l`�1�i�H`���:�%�\]y��y��Ƭ����A��,��m����S�i;�k�8��|��6�0��g�E/�ptzy�#���72��CDY��Kwad�\;���Qo$c����o���������ז4�z�jY�@�g$���"DP?o\/���b�;�i�$��ywŌ 8C��t֦v+�X��]��9,�4�ї"�ZL����?��F����i�(x�9u�[􍏪�:X^չv�'��5^Ne�<xb,�����R{ƋE�yr���m�"�W%��� �\����)[˷UkN�nxa��pz}qp��"s�cE�jV{��Q6������\ٙW���Q��M� ���wi�^���!V_��:���F����a��J��)������%}���\h�^�TR���_5*�n�K{��q־�;��|k���a��hH i�o�
&�U����DR�����i!�|0|>D��>}�=�i��Y;�:;��tk�	��P����'V��&v�c��D����i�
(�������D�KM#���	NJ��Q hup�����I�c䄐�tc�<� t�0�"mNI ��2P�Uh#0���$��Iѐz���PAi��U`���~E�$c�OJT���p��XXa���;�)�� ��8�U���xk{�es##�cY��&���)�]zs�!ԥ����J�<�o��V����8K�p��u�3q��+a5W�`bԝ����;'{x�݁�S�<��˩���S㢋��mh�[�p<����,�� ���E��T�t�[����h�h�{c�x�N�]�G�*�=$�5�*�=p���(%��3��ϧ�[��@�_ �_�W{'6T ,�6?A��3���6[�J�قs�"!�$ǂ�7�D��|<�ڣ+^W��[��n�yŨL����p�h����T�N�v�Uص8��d/fn�������0����|��x�U�����:< YaQ�rJ�%!(ɁF�R�%��ǌQ�5�0���7c�[�b���kMa ��'1 �ଌ-��=yA�X)ۆYW����5���N����M���=Ζ��/���^�}�?��n	��;�W�N�EŁ%ih�����A�?�	��vĝ����sk�,�V=�RkY��*lW���/�[�h��Z�._#��b���|�����%T��9���Pg��~h���U�P���JCv�� u^�JD7�2�������'��� �<Ț�_�^���<䖐�T���C��һ!��i���'�E�+8y*N�!^�n��rCo.8�S��jj��ۡ� ��y��C�а>p��a��j�\sp�:kBlsCh�)�񷤆�j9Te�b��a\�@�� `�cN���Q�����m����C���R���'�q��jqT��[�5����}�����%�}.4����W��܇a_��F�ÏS�E#v�4�$��2
��\<�vt�����2�mNy�����$�N��
�ۑnE��H�3���
��f4��'h���(fJmlqS��"4t���ʼ��}'+����E��2�?�}F:�+PKƒWI�Ur�\*�*�&�4��Iy��!��o�t+L�5�&
������M�B��=�5y��ĩ=k�xD�����.�#&�c���"DXiVtH���Y�&l�Ա�
w�c?1���	w�� I��t�~���g�>���a����C�ik�
�f��!��J*<ם"k�y�Vg�i��%s��25��<�Q̇t#'��in���[�t��լb��)�����˕TJo���9/u�"���ZGw�VnP)=�ѐFM9b�ǸVKҒ��v�$��E�5+� � ��������Rܸ�P�=����AC3���-�Kƛ����r�?[�lVj۴�6��d�߮��A���J��,��C�>��RG��L�����J�w=��G�<ۡU\���Ŝ�M>e���I{F� 0���:��_��AGWP��{��yj��f�Rf����-�[@�^N��t��%4�7��|��H��t�0��V�'�:�x�(�ΐ���qH�oó3�4K�����|'kGC$�X��t�']y�B �b�h:$|�	T�v�.���E�=v� ��Rp|nB�#�3�����џ���?ժ>�[i�������2�0&�]��p�v�a��|��+[���p��ٹ_�bׇ����z<x��Ը��.�"�%P��l����?���� 6`��R�W��Qw?KM�� 	�q��ֱG5ːw֙�&���Ȣ᪷�k�
Qm�S�ˍ,��D<�;B�O��`�-��������|�]���Uɓtތ�5g@\�y3��?��O��Pvh�C�|b�m�� H�����3�t���0��E�"	��T��<Ӿ����!2����X�E<�h'6�M�ESd!��1=aY0����q�i���PW�R���%���t+է���@)���2�ͼ����OBj'�%H��k"��z��UGznD���E`��;6�\&#����l�)�g6�_�^)*i�����"bu�PC �(�6�I��9[��