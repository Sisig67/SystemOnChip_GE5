��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQH�x�U�'�'D�~�U�:�Jvx6�v�h%i8\��^EFP�еb�w-"N�uc�v����aL�r���n0n;����#y�z��Y�ZT��ϻDn��*��ܒ\��F2�c�W+n�{��_~j�sm9��h��F���i�#�OOpf�h<�b�$,גW�E�(R�#VL}�o-�8Sz�\�VX�l8�r�H����3ۆv�����a����\�ԉ��#������Н�����!��\&��_�Q��B��8)�q�VƄ���6���4y$��7��5�a6M~�Ϟ��6<���vvĂ�3�����-)�7�� ��5ác>+����g�+��w�zׄk����_���:��t�vmm,�����n�fX��ņZ�4�r!I�je�E���N���2)��efb��98/��`k]]��Hx����T���y0 IL�/#�I�z��2�8X�5궄�-_*���^�^i�>_��$i�8��f-���V�3��U΁���k�*/�����%�܆�h��%�~ݯ�Y�}�z��X@�q�O	�w�Ԉ_� ؤ�Q���=5�����c{�/ޯ39����H�y�R����,����̀�e~������<�ܚ8�K$Ǡ���BL)�socX�BWk�?E����v���ǌ&��K��*j�z!~VB��%�v0�j�/:�t�V�64��c�q?껹��Q-�X���e���=�=+��ы�e�&���l�G;n�"�+�XD�>c��)Wm�4ɋ�IP^O��Xiز��Aݸ/ 22��a%�y�:! �M�z��Z3 w"�Hxأ�:���K��\��G��Fj!�YF���w��w��O�a�j�����f���c%>~d8H���BK��6U�8�Q�G!�l���dFE�k�!�c_�{���Xxa�ߙ w��-��"���MX�)>(c�L6�`?r�'iy��p��l������^ͧ�s��A�Ew�m�ׯz(F�����:	�>�3��)1~Qpn+ZM�<Ґ�ߞ��hW0�q�Ӱ�T�VU����2i<��Vein^��x� ��2Z:���T)A�%��M5��yX�����y�'j��;�^c.��^.���c�L�S�:`��`�Z�;~R4xxAꃡ�#�z���(�epK%5e��O�H��ΟE@��@�ɴ2��~Kk�ъ&�j����ƣ0��z4�X�5e�x&ÀF������	�����]қ}^fFo��q�S"2��(����%���ʒh�tn�D?�`\�!;�����3��ܡ�p�3��O�*��2g�ʍ�bk��yE�ے�<�|�韌���8FM���P�aD�f�K2'��Gl�0"zh�Y�`|��9l=�p��*|��i���V5Y��&f T��'5%mG+�Rཫ��[|GK�q���;�9\0�<�1Z�m��>,���+KpO�8?�21�ePθ��I�O�J��;¡km�1T���J:���Im�)����
����A��W�S޷��9��}�dE8-���v_���1;-h:9�*]G®" Po����5��:H&�q�X���c��?����b�o	ˑĹ�$Y��rz	n�f!"�.�^�Dt5c:�s$��ÿ�� �C�
;`b�%`��(C�,;\iy��թ耣F���b�盢�ǸN�q�����PIWۗ����G�Rwt�C�N1{�a���hJ�������f�$ĳ;M���'�[-�_ ����#��;?�R�ΐ��fJ3:���&���2���)���iG8.���4�&���:�]3�ǁN\yT�4YulnT���]�B�s� S)k��'x�~��%��uoK�[�/��Hgz��Z���Xr~T�"3����r�R�2W�b����ǜAڟ�`�Sw�l�,y�����rM��˄�Y'�p:���UK5�~��৊�V,�Xu��J��L}�<ܖ˞U��4HQIdA�5|t����E	hzZa-&}咢�k�d�wb�O��zxF#k��N���� �R����u���)�W�I�m��5�i�}�O߬��~�|��yv'�BO�~��i� AI�T҂�$g����Hn��nE���釘�K�`P�AK�?����M���ذ��E�ĭ�r�g_v� +Ռ��s�w|*�9��ͱ���)��?��]f�΂�jr�+�B�������;bhE�\:�ܥ�8�� ��hy����BH%zfѾp�1��w�ߪ�����)B��׶�Ly ��Q]�;�n��Ү��u?�u��tX����lc�!�����'�A���V�Hc,R�t��{Bn�I:`{��um���������ko�{}�߻}��+����v�����s�D��F���:tw��O oyҴ��ֵV��o�����E�[u�7�\4*=?hV1"����v.��g�6�mѵ�x^��2G�x�����/�&�=�	|j��,����\Ru�A����-i?��x����N��]��J@,�����4� j��@�
�#x�ی��a���}�A�F^���hDk����fI��[���`*㢹����y�38V_�Ҙ�:��#��0a�w<�r���^��?��.V"����]��N�h�W�s�d'����L�v�Y�� v����	��c�<n*��6�{���aߑOF�p���o/���vD9�;Q�%��MR9#�T�{��śd�Y�2$��]^����1vB� ��vM��)(MV�\.�<�dd`	q�5�C�n���k,H|�9�{��+���o��KX�5�5A�����3<a�#�о�߷����:L��-�I0%|�&�p����*�F����*4��4�W �����4?K+�S��^�1
�l�T��o7��]�;ܿ܍\`�,"`���y����{-�&��OW��4���f�t�q������(MU���7�-�p��I(�⬂��c�+��Άt�X�$�����t��1����� 	�Eu��H�K,YβW�3��}gI�҄x�Pu$Ye%�a�^��;�m��0ciJ��*?Xl=��5�d�k�H��s,˦�J�)�B�{�p�bV�Qp�;��z1F��d�b
�ق���75�~=�>��� �9wZV�S[	�r{��9SkUl���s�V. ���YJ��-אu�K���DF
�]]��j���6�%Чwɤf<�%��H�i��l>pR��67��H.M���n7��c	�h�g(��W�G��=��z��3���/J��+P�;��!Z�~�=��!�D%�]ޛN����y�7����{<�PiӪ�FM�+�&��!��z��E�n\J&Z�L��'��Y�������|Y���e��M������e�G_{PP偒�����ì�����(%#{���(�IZ\o ��lc|����g/s�W�D@��� 6���O4����'|�?�q4��z�aGԌ�zq�F��۬�iMCB��7�~�Q���ek����g{�&3��d�� 
����,���cc��:��t7��وMAo)�x�{d�D���q#��=&�a�u��اKri�~ڍ���k:������������7s�&��g&<Y#�X#
��=0��~J�8פ�w��w"�����|�����3s���3�|�
����OTx`$�bw}~�J�Z���Q#�M&���^ܑM$�D3khT�*6s_QiB�"Uk�����voE�}��u�,}?�|�̮\>�ĊG�����~ʣ��V�^M���S�	�#;���]=��=�1�+��;��Y�s,�Yԑ��@	�vD�ȆB����q3)V;���t6���zF��|qQ[�rJ��Af�mjZ2�֎՜���o�Fs�g���7D�舜$��y]��/R���?8�ҍ��L���=r�����r��
Da��\3K��9&{,%����W9��%3#+m�>qx�6ُ[[��u8�( xx�-�"1h�Y��E�:�;-, C)��-=�a��d�������+^1w�=$x�x�8��c�*�Қ٭6�p�떵=%G�yJG?�T	�2 ����x����Sg<h���>z��k�n ���.I�a���o��y*_v���S�f'����4-�N�U�@����b�<��V�����([����!#D �\���,�Sd���y~
W���c,b��G����
�sk��a�}߳u�X	�$���8џUSL�Ow��\i�'����Z��2��0[�d��HV��j�!h
���l5A����(u��l	+�`�I�B�T^N�:Y�,H�$�:�R?�5蠥MOO�5$�pP�+w�oD���m���z&H�$����C<{_��t�D�� �`���3�\�ig̔w4C���� �!/cÀ�g�z�:^�h�m71����j�P��#���k����d��e,���bO 2U��q�IF���!���o��L�v���lo�5�0�m�Ŵ���meR��X�` �a�x�ZY�Lf�����t�q��P>*|���P���L?�i0_0B�Ӣ���T�ꩤ�[p.�y���1�1>������� ���ʈ�тH9�9ڊ��T`?��aq慘e�&�]�U��Q�-�
aQW\X Y�+���r$XUE�
2A�����.w��?���@�jPK����������pޠ	�����='
��Q,;~G�+����ȥU�!	.oʧ�����3�÷�A��4S�����W��Wӓ�+ʯ��/}��{�假1ݚ�~@<U˓9��}�?jɜwLo�2��5/*D�I�/lˀ'�I@2�������L�Z%.'<J�#��a���s����j�=�H�dIDu�t�$��u��xA=~-V����.(�j]]׮�#��3���,�A��6z9E%�7�8��ӯФ������7�'(�R�|Ӊ_9W�T�t�c��	�7*~p����'��EV��OىDD���-��=�,�Q��(Ϛ�.��Es;*M�t�!���֍(�']2��BQ��b2ܱ�a��pg��%�S��'���pa��(��{�Fc)y� ��=ğ�zNP����'�'�M�ኰ%��m�3� �	�8�W|��M���h�eA��ߦ�=_�\��9�@�v)4�������Qs �/��E׋q�� 4�����5[�������\IӬAaF6������j��?"�3��t
�j��s���H��K�����5�6����Qo�,��Hd�	�*_��i?����ۈ�bڧ�Ƿ;����'Wr�c-�Y�!{��`�q�1f�����GG϶�Uq5�M�����1<<=�n�\G���S���.�goM�DkO�,U��u�IϿsY��dF8A�D���8Ǻ�Q�^Pa@z���V瀥ʍ�|}W�?!W�󢰍�2!7$7�<2JF&��(�tW�y!/�^oUs���Ꮁ��-6}o@�-��v�����x��a:�m�9N�c����������9v�J�N�f�t�Ŀ-���\��=R]S����,?|�������d�ڍ���Ĩ�ԋň[И�I�W�l�!�� ��OHi2�Y�M�r���y'�2�(�#�;R��#b����:C7 9��Z�{�Pg!	���͋�4����F�=��q�v��K�_h�n�Ņ�nߺ�f��Gō��P���M
[����'t���oIW���w��hzG��0]i��D�/Ғ�X�{��s�v�f�؇���t}�-6&��o�_�nH��x��+wy�Ty����e�Y#�8�t��lM�FF#�*�7^�p$M~vn��p!iԀo3wDcR