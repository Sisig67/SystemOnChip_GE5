pll2_inst : pll2 PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
