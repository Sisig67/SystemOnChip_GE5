��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���|���Y��w�粒8k�о<�Y?����tz��z�I�y�ok� ���j9W����x�S	]�`����SC!��J�ā��V���� �����1W$ ��r�5��p�?�|�����G�����H��Fgõq/M�F���Q�B?O���������bIe�seaq�p��*G��xFi�Z|U��%��if�O���+P�pt=+ ���z"����U�K�l�i��$u�)P�,����`�2pPNk�����|������?-�J��Q�f��X�����ߊ|��#ǉ�Q���G�w�j��D4���h�A��L[�I�a�A����tZ�+=�H��=�n��~����8s,t&���eo�<Б���W�S|mIw+-�������Ym�sF{�WIz��Bc`�Q���b?<�Ð��R�=N�@�Q$�����=�i��*�M��!ޗ��p�^N��}��L�[d��OF��}�G(3!$`��9�s��f#D�v�.�pw�.����U���Be��R$�	�˻�~Et
��I:��X��#צ��v�tg�h\�ɞ�I���\��v@�_�uM�s���·[��e���l���^�Zk��Å�$�V��΄�^��N��X+7��#�&B���������D*4=�5Rg�����{H�<�6/����!>���NR����L��u���jd�"S��i>���(c�)~��7S���	@>�¢��ieQHN�:��n>3*��N4r4�ɽ������x���)i/I�a�8Vz~bRKQ�3,��~��`z�*�V8`ې�a{㨴c��[�6)���9�q�J��=n' �˚(s{��4�9�"���A9L��)"9�̤���#�������n�����XK|Z%SJ�!4�4�P�[Sh܍ϴ0 _�F�<]Ҏ��P=Ü�"N��4�g2ݎ�$O�b��0=��9��Π����-��c���8��!k
�����Ŝ�=c��3���������'b�u�(F�G��5�hk 
;��;�m�%u�v�IT�q��N�F�XK��f���Ս���N�����}
���ma��<�0#��u�r���8s`�[=	Rw:�ħ�x�F��mg� �*7�4����_,*��_�.c�/X���o|����US,���#@��Y��跳�\-�}��2հ�?�?�n�c�JEq��<]�� ���1%�b�-s��|�-�S�_��v0��7Ma�)4 )J7`�7!�z8����J{	oHq� ',|-#�:�G�x����)ٽ�Œh�D���!ܨ&�ǭ�^x�����1���M
R�)$�����%Lr�DR����i�왐��5��g@w3Ѕ�O��r�`�c��O�S��"�4���Vm6�Myކ�VX&]�]��t��B.Q����%il~���D��M�P��p+ĕ ���9:St<ȯ��S����>2�@z���Av�}��Փy�O=�)��k=�:���� �O^Wvt]��[0kn}彡M6�Q�����2�1����+xe�8n�ج�{V����.46�9���uj�������vcБ���f�\��UN�b���z�M��{��Y�
˼ԍ�8z�|��z��f۔��o3f0QJ_<d���1Mɜw�r^��j2Fy��8Qmʚ�cM�i��]����QSՆ����fP.5�R|��L��iY�H��\ =�7
v�h{?S����q�g��sAT����y5��� �ε��s2���
vE�'��ht�}~�eğ2���K�^�7y1D��D�NDԐ�LW�� wD��ހ� ����6U
f���;��y�S���8��a��.wGoQ���I�!ǲ�\=ҒxH?i��U-.t�ԕ
�Tp����f?�5Rk��?Z�s$�ly�� ��E�&�9E��Oq��ZH'�\?q��wU�{�E�>�&�C[zq<x��s��S�9g���j8T�.Kq� �(M�!K���mF��NX�I���!o�=[*B5<6뛪͵:F]�Z���Ѕ4��0�
.�BaI�+,��Ll��q��gT�o�Ҫ~/���I[Y��U՘�`��Y:W��/Њ8�&�À`�V������f~��d�uuY��/.?�Y�W��#�R��/Z��#6���;+"c7'd bM�9~���.xb<�\U�_� ��I_��y�z7A�i�����{L�WJR��-	��}�g�J����rȑd���[ ��h�><F�ڈ��~Z�4���עlWSo���4Շ�ǩ�	I���%����Y��R�`�̷�4Y�?���4��f|��A��b	��W��jHY���o���Ǣ���o_)n!���&�I0�A���w�yrG	�#�^�N���A1}�%��[T��x�min�ɑq�q+L횼2$y#4����U�����ݝ�O�`���V�b��1�����ϖF�s u*���-��2A�^#ro-EjPy�rz�,�*ki�y�'�H��-�S�e�ը�4�h����RX^�n�i�R뀩��e�iNX"96���i1��`ś��]F��+�}���^J��o��fL��B��,�a �j&27��`��>�V|w{����2 ������c����VȨ�p*GUC����k�g�_YQ?�YO%4��1	\�r1x�����:1�)d��h�������0OPٸo�w!�Ͼ���1����៴o�@e޵�R�7�R֣U-3��Q2�휑7Wk�Ư�;���w��,E�Q�E���ck�K�x,�H'a�9���9S����W���o���:�qX��
v�H��8,6?��~�&W��q6�
US�Wh�:�3J?��g�,�^:��h�#BT�����}3�n�u@�O�Sl[�,�+��7����unYЀ�VL㻲8|����B�J7��a�Z/z2����	��e�g5�lg�����I� �`�G/�B-ϭB� I4j���RU�Y=�"��`��� �h�>��x!��S�h�>#��f�e�\?�:'�ј�}��B�Y�'8!d:�(a�<�j�L�(H�W����D~y7���S���[/f�JԆS8��V��`:|y>���1�x(V�9� '�%�ft	گ"$�$a�z��h�g:a~��d�m�3����˱�w�oF�tJ����x�%�Hyo��:�)�	,D� c@��1:2�R�Չ�1�E��ڪ4��a�V��2Px�"O�Ե�@�C��<�z���8���GfˠC��},����"��R�W*a0e�,�o]����=L���f��I}B�9"DP�G��{S){�׾�}J҈�S��F^m�+|y�����R<�[	P��uhI��޾��.A��!��v�^��a��󼇠 \���Ew�gj�)�A���l$����aD������m޲6��т.�@�����J��c�=��
>�<�bk#*C����5�~������X����[�gF@����x��Y��Ch��N/V!��>_z�B ��UcÈ�A���)GS�9�ǧJn�	����e=|I��ީ�H�#�3���f�T��3�((�����+&�UU��R`�����~����?���0k��$�Q�笯��c�b!���.I�fxύK|%�e�#D�s��Ω	�^z�ȝ�!d}���b��,>O8o��Q�Gb����bxr�
9��N�V���7֣�OD��|��>'4�cpͲ�\8�@���aY�zl�M�-�|�[��Z��{m-�k8^�Pu�G$�h�@�h��P�-Z�-���7�m9�:��Z|�\�:k�i��>d9k?�ɉcT`Ͷ�}"&�i��	��v�o����<hd�a�E�t1L����^錤'��Q�'
E
�~����sf$���=S{�{�О7�Wd��@����qX����<E~���$���t�C��d�ʹ����O�w`ҟ~M��E�X��?��5�bERL�/��ˣ��7W[�Z1�6�Dl���2�Y���v7P��67�����*���+���#N�Azn�H*�UO�:��c�xy��w�m�:�]3��c%g��rU�zecQ��8�c���W�\g�C��n�m��fw�_��[黹#��O�MgO��I�/���YZ� �,H4PD��-dU=$�����P���9k�/�Ӡ�C���3����l�1���zo�Q��nA";l	�/���X�����6Bl�T��;C=[�C�0�0�c�tU��?���뤽�Wt[%+��UD/幅�|���auoxP#�����?y��-��βB *
���N�H�Q�
W|������X�&�N[�����X�gB��d�Y��9��϶+��K�Ӵ�����*�![cf�b�{�ŏt<�˱>�,�Mw^��%�!r��7�u��28�]Mv�۶Π[w��{��D�bW~=:]�]����X���B�����+G��m���z�=��͆��b.7�ra^@��9���6��g��D��qNk�Η�.���*���v��/����b���D����4��XXy�b��I[p�o�p���Tt��sg�M+��?�mPQ������P�9��0��ָr�O3��pJU�u�#g�h��{�,��cw������Wx���_m�M�~҄�E@l�S!�B��䓿5Z>!��d�q��&���~��p1�ӥ�����n��Ѫx����Vs��4r���NѡhmH�ɋTSU�*Kԟ�A/�s���U���s��}�
/��Y1�W��	�	�9�s'-��_�r�w�I\�{�����&8ܫ�d7[��\K���d�S�G�
��59.�@�y��������Xh}�!�g����_e>*�ؤ# ����NA�+����n#��߀�*�Xr�x�u�g�0'[|�2K�iC�uR���TVO�G��-L�{��mW2%z�� 1z�q�7V�@I��l��/x��[VA����k�T��>b_�K����~d^ٙ]��w�ٟ���#���.�߉���t�_�F.�TgN�p�Bs_E��H�xOۉY$�P�p�����LW�Ȱ���	��������JN�w�R�
�"9��o'����4ykG��ޯw������Y���S���CI��W����]�.(�A�mR��c�IҸ$M,ؐ�e��}�'+��i4H����}e��92�jt	��*$�_�zwKm0������d�2��������9��$���"59��^�۬�J�W�m�^+���m~P͖�-вȎI��(�������G���{�a+]<]wg;6�9��{�'�$�^\LWB
���+����<��.v�$D�\{!3�0%������2PW���`��Ҿ��x;� ��` ;�s(X�yN�uV�U��=,�a��}�iz6�[9U�"�]]���4���H��"��κͩ`�����i���-ݟ�"f<�9�-=�Tl�#m�,�5�,���ҟ�T(�5z�8���a��Ƕ�:����7 �+%C�Շ�