��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����� ���Z��q�N���B{��!$���W�f�Є��@>�e<�e�����Yk(!_GN�ν(�	::�b�^�'?-a�Rɜ��Lm޴m���Rt��z�U�7�&��0}=H��z��Iض�����s��LWqdJ"ܳ5r|�&�E���mēm���͓>��� W��E7P]��rz�aTq1II��|,��N(#y�6������Mp�~臍8]�o��:*ۧ���}q#��=���x��ݜ�)v��a���Z)��]�g9m�j+2�G#P�5":uѮ'`230Ґ��¹����>�����fϧW�Nz�����Qw�����/���5{J4;,�}�0��0��z����v�,���ʮf]�ϼ�狘_+*�v&�g��%�M�����;G�F��,��O��cPK/+1����ƞ�6,�4:�I������z��1�S�
�=�^l��),tg��<�Jg�����������Dʅ(�G-�7��&�hTRq:�n���ښ����+��C�	�ԩoؐ�N��8h�$Q��`V���{\u������*�����O�M�X)�-���8���a�Oi���Al ��d�ţ�!����Ŗ�����B�0���{�a9]�oͦD�lՍ2�s��j��1��hS/���H����u퇤j�-BS�Y�を��F�GN�~_��ͺ+r�Jy�k�[�·W���z	Nj�c9Q���[�"�E;};F��{����͕ B�~z�Sm{U"��� �=X�[`LF�.2����BP�_`��3
-����-k���&�:C�;�"���ɰ�b�ŷ��5�Y|i��0£����{��A�2� Lߖ���QI/N�rԈ���Y���G��,Ģ[g�N{��XZ����K�="�}W��(]6���c¸-�!?j4�%�j��Ʋh�cB螓���o��C��q8�����A�Ը��@H�2�j����λÆwc▻�r;�Z�	f-S�c*3��~So�R[��J^V��ӡ����gJ�[�Pz|� ��P<�yD�l�g�k��X�V�)�8�w��U���9�:.�I2��ư�IM�U�?�T�☡����� ��Xm(.�]�'g�e�I���I|S]{�۱���(�{��^4�9�f댂��P#�B�K�yAe��E�!oa;5�/V�e�t���D�bv��X<��NӮ�wh�P��^Q�b�߲�D�qp.��m�v�q�ͯ:��_��~�e .M`)dq* �M�PG��A3���)�,�0_�	�`����M�:�-I4��*�qo_�+�x���w,���d~{h�uT�<K��J炡m��^��G9dcm��	[�i�S6���a��������|�� ë%?���~��� #�ޘ�K��?0+�_#�2u�Iq�#U�;�+�XH�X�)���!j&�-�L�<Rx��>e��O���h��$�6Q��jlir��н����Ӂ@v`�<�Bd��Ae��_.:���~B+��y2�b�|�` ?�����ZD���3u����;nʁ.H��Mi[6"�m.38ª���`߾1I�!���ڔ�����O԰��=��%g%d
{�U~�6Ji�D�9OQ�j�+ ܮ�w��b{�Ī__��h�E��{���py�)�J����΋QBN�Mv���Bh�"�� 15?eT&K�@�@��X�efDR���Y�`�f�"�ȡK�5Χ��bd�-�n~�����t��%���g�zq��wٝ/�{����Oc� ����M���o�9%�1��j����B�&�������:`o����,"5�"��.2h�� �����nж֞���� <����y���qɗ�D��e6�y�r./]1�h<�[���*�GTXHBu}Z�m�-�P���n�(u��{?�ʍd�g�5�5�{��w$�4���`�����N�a<����vҚe�y@�#F���� ����JNxg�����K�2�v5j���bI����V=��3��D"����y�g�p�;�%1[�r8d�P� �3#W5F���� 4h'�;�^9��7�Є��XN��>Q��W�D�.�Է}lo_hw��2(�yܜrA���;�g�L� ��[�.�Ш��]��r	��&�B0�=_��pz���9�f�P����+k��P�L�ԯ���n��:�ʃ汙�����A�B3ͣb5����5�M�fZ>6�͙z���0~�K�m�dĸ�d%]��������2���*Gi�����D�壌Y 24�E�[�v�pKkO�@���y�M�;�P�= �`E���]��Ȇ�9������k�H�4?��T�?�=���/d�G�fz?��2��2۪�xpK_�u��,&w��K ���y'�%���U�,��?�D�K�tMf�?f�$G�JE�n6���#�2Ŝζӓ�G)�y'p����G����q�sދ�'��f���*{����!兙Z���ւ��g�h�D����#�q���"ap��
�$�9�E&���V�e��/ �-���e8�W��(�;!ʠ㜶��[93*U�\�t�#�I���<�{g}�+:��[)=��nB��c�b�[�3EH.���J���%�x�L��C�Y^L7��6�y�~�v�d��p�_���-zO��*!���`�s�V��Wj����-�s�V����"�"F'7�d���Q��fl�1���v��|2'�r��a��ά��Q�8$z��}:��h��\��`(Y��:wOx�'�p�؈y��Żk����� 8b�;�&!!�����ze\�%����Z�(oJ�-����U;T��ٟhC�#�|�o7�&�%b���Eԧ�Ʊ���euzH�UygX�6�n���Uu�Jrm��� ��0#�)��5S��D̵�B�
�ג��zG�X��q���|��i\�H:�%�6g�!4!ۜ۔^Sj���LNu����ſ79Y	]V`f���+�>f�2Ϥ&;�m���q4Fs�v$`4릻zE�c$)N��b� ��u"��K���O:��4(.��3}ʵ1�{9]7�q]�8R���t��+&�������YްF�{���7Z�!o����/�
}§�2.R�7xwKX�S��ߛ�����DP2�*V�h<Ģ�DD��!l� GֺG�%��E�����"Tɻ �%����'ڧNww�s��H��t��`c@�1��\��U�0�����6M�\�Xeh��>@V�b���f����ي�#oB��/��I�K��0y��m���ѵFh�e�3�cjرn�W�xV�By2U&]Z�s���LŌ��P�3iI�����WU/~I ����\��-������)�-�4�@/��sW~��Z��]������tt�S5�����h��d�,�����.3���Uopx�%�'�X�j$�l*�1���_X��~��&s#�W翢�O9t�0�h����К͍���5�I%�Vr]�m�[Vߗc���믧ݶ�1�C��������F$�t����/�-UMW!D3ǅ3��5MEn#��.v��'v(�I��i7J/�1�&`-�L���i�a�yK� Y�'�D��o��N���|�b�{La>�Mq)���\�o�gȴ�č�|\�6��@J��7_�� )/��ya�x?{��2������T�uj��d	\J�=�d���E��	3�����8,j���;�D�A��4O�P ~R	����>-����n������M���V1������Z��q��[�ZZ��L��{����#(���KN%5s��ҟ�=]�=,􎶮��/��Aق#�p��l�[L�[{/Yc�,�h�r�J/ls���Qr��[Wm�����=߄�H����&\S���� 
�ݽ0��U�!��!�G�`��B�+'�4���W޷�"��#!�X��G�����{��SV���?"e��o�|��v�z�̅�B��@��s���kb�|�BB.�����M�5�֟?�P�f���i����� �8V�5=o'��ܷ�����q
��Ȁ�˵$Ց��#1rU�5�MsuJ��v��12��h-�}b�8 �x#PXF�9	�JT���&�[HѢ�Ѕ�'f����ϲLڞ�3t5k�����Ս��{±�� �O����l�+�A뛔<jD_'��o�����H6�&��f�Pi��~y[��v3i�y��~B������(}P��f{��X^����j:�̄����햫�I����5#%�uM�ŏ/a8.~��{��M!�#�[�)D�5K۬J��q��Бk)ԫ�^������n�#	ͯ���
^�����}��ʒ���l��R C�T�c@��뮍�ʐ�q:�=�H�����X�����"*e����o�;����M�ۣ�P8Q�d�xdǤŚj0F��Q-gNT��C�ɯ���D`��m�Χ�y���x��2A?hhp���"�G��P�1� m<(�A������p gFu)y��s�7Q���2�+RxL�@mAD��C��.+|�9�����[Ȑ��q��Nz�X3�YE�:�G�|f�p���/��,�(��
1�p;��y��X��?
A(`Ժ�'X'MF�?r�u���E���#�yD����ۧi�f�D�g���K'.�F����f��>/�kS]������l�Z�W*��i�m*��A���o��	c�/TA�X5��T�ߢ�qn���[3n�^���{�Z6'���һ-�`�����ٖʺ��EOX
�cKH�
�l�w� ��(�,�@�/?*팉Z��+�oifS�)�;���)�b_��������R�����E$Ɵ$%����6�8��uC�n\�^��q�����巚F�U��Ϩ:�X^Zm�]Ð6$	��G�G���	�A�ا������Z���W�}�S��luD� Fk!W7�r)�&914��H��d���.
RfK�Q�t�*h�$�_�di����qtm��N�zd!�~��ñ�sZޏ.��;�c��*g�+{�:5�E��u��?��=ˣ'a�wG����RV�E�ܔFT��;�Y�u���9�{.�a�|�hT����{]��W	[�](`�$�`��E���oL`e�P?�X����[�w^#j��+�w�@�����ֆG�<�Ѣ͟sB�y\�1�Rl΂PL�/31��m��#�����Y|��oL�-�q,;�ſO�&��0��Q��RM��Zq��ҐH���;Z�4�Q�0QX^�6g��V�����n�D�m�� 6����0!�h~6;�zG�Z,�1����b�����;T�`+�9N����¸�U�s�Fp���ȣ��h(����ٞ<�-w9����c�М�]���n�kS��Vc٦��n�I�LWo�kA�
����24��}C��p�
�cV�m*]`oY�^�` ٓ:t��C�o�i���0�,!^��!������H�ӛ	�d��I�Հ�V_����������CW'�F��Qй@d83�rϡ���uD���8����IFAܖ$WOq"R����T�A�1_4��6�_GP���>9+Cu��i��)^}�C���E2�مv��M`��)�~֬�!q$��"���n��8^�B^|���f����
�G�I����v� ��p�@^(�Zt37��5���wq�G'.G�Y3�\�d�c�Z��!+���)��e���������Y �BZ����V��P�l���L�0Tv(��J3����v?�c��P�	ckk�$���:��}
[��eK>��6�io%��(�� �����.q�9�a��p�� �"iՁ:�N����[q_�Z�Z��W�����#w@�q����%����V8�{
��Xf���Ɍ�y*+oNI[���X����J��k]T�y��ő�����$%w�i�+b���s�s��$`\�v�����q�a(�];G��~5@'BK_��
6SG��?Ym�PZ��nXl%�2"���ݏ/^a��EZ�����< +h_Kl��:u+�^R2s*�NM��KI��$�,ݔ;ޭUYAE��b����p�R�B�3TKXI�Tfz�,� e�I~�Jn��V.�����P��%&t�_�%Ӯ�Z3-��<a
�!���)Eԇ;�h��M��MNb���f_o��\�q?ܠ��}�|�7�i�;�@QS.�?* �.3��!��l��ر+?	����X	;�g֠�9 <le'(c[��AU~T�Y��1d�;Qu}lU�����@�y<j[����X�.,0Ti<S姏v���>�9�W1RK6W��+�յ{�<�6rL�z��/�3I��B*L桡���@ط3�
��uMF�<�'%R��v�Puz1��_5N���*�im�ɕ½3��lR���+W�2ڰ�A�@���Z���b:U��9�#��6c_P�2�+,�`��ܯX5��sUM-a�-��j��a����	�0�u�l�SZ=Y��Y�F�e$�[aH&)	�ݜQ�8\�
s�hbx���o�������҆�����V����~�2��y*q�:d:�A��@���<lf�*��0���<`��H�B"}�|Ý�	@����x۞�S;���F�	��Z8e����� �F�=���?�]{H�*���E1�C�
���}=���ĭ;��sA�?`{$"�<:g��s>%����<H���I�i��!S�3c�8tG��E�ݺ|Z5��x�ݑ�Ne�^��=�rF?:i�����'jQ��k)�2�	�A����'c_�6�L���\?l�q�AB�Z���mٍb��w.D���b��4S�|zꀵ��-Qu2�=R��J[;�!A���+�T����d��A���c�	3T>�E� 4H�����Y��Q�U��\vD�{�����wX���~2|�ѻ)�2������I��K����x���~.�C���5�y<+�䒁*�'���ӌ��CM��b���K��*�M��\��E�`�U7$d~����D}BF�0�?!�¤	,N�OevH"���Tut5/C��2���b���p$�7�����$5M���+�����5�)+,���ul���+�Ɉ�k�4<���;����l5sk��7�)60r����~�?$�wҍ`΅���n��S�u��4����h?��$gL�[����O6������o��p�t�o�n3|� �M�N,��,�c�2<�ХV���m�qp)ņY��*�v�����񂝆�ǄKǻ���'2d��tE�z[�a������V��k������!%�-�agA���&߀\K4XV6�|F|��r�[{
�=�U�I��wxp#��({�[Ϗ�x�3��}��{TAf'��~`�$������~�Ӓl��r��g+c��w�+��ٙ�ŕ;a���;�\��j;6�(&��@]&3��x��� �P��%8#�v�чɏ�2/Ԍ��㡩��x(��_�q�^$_���'WY�P��X��
坯�j�����̫y��c�r�,���A.�]=�^;�#�7�E	�nD�EC��6K��1�����f5��
x��#��_�J������]��~)��w����̛ {2���5��)m��)�y�n���Y�,Lw�\A���]��.��ݨPb�oI��tu�yh�Z��^� �A��\�����3��YL�
B�������UUGw�w_�w�(HOC|�M��p�0[�l؋]3���"#ht��*���3���5FT�O}�7��CYB����3̅ٿp�sX����A�ou��؊�ȡ�J��f�R͓��5�y�NffR�?���da��d�Qκ��F(���$dњ����7�z�����^ϣ��g+�-Y"h��g%�Q�B'J���9D��y�+~���Ӎ��r��Ũ$q��I؊�j+W]�~�P�U���w�O��ۙp^���5F�'d2[]	}Ų}��L�6�1�S�f>+��k�$i��ī٫'�V�VzMQ��Z5�=���8|����S��i5e�r�'��>��)�~
�z���цV9y���y悰�J�m���1r�W���������%�)�?&XA��Ń�VM��IV���&S($�t�����*��Ǳ�)�P��	4�yT}�H`�u����t{)�
�p�+�_����iڣ҉,eƃ�'������U���AT h��q��p\�2/F��y�ʬॆ�X0[-݃��_�T����i�{�n��;��3� w��ާ��w�V6O���BY���v����d���n�(I�W�P%
}�����w�Q_V�@����u>��'�����H���@�*���������#�t�(tG�����+;h�k��씾�74�v-5\��M,��Z���a��37m��˫D�4&
��
�yD��D{��-6_�[[��H�Z���^���^������X���p��{���>8݈��\&6J�:�������V4�OU��,�W,�v۱>�3�v�ҍ��;�¢6�6���)$��h�����պ�!4Ӧ����BA{����
���(4iC1�8r����A��9{ֽo�+����bP[m�<���
��g���0�?3�"��۽[��>��62�m�u6>���r�!^���h��:�	��3-	�L�x��r���_G��v���S����ړ�%u?�Rd8���|���Ԗ�&c�4R���'�ym\,	^�,4��{���U�D�"6�'�h�r.>�pi�B����ZzL�H6�r`r㺣�[��� @�f�Zٌ��뽎V��1A5�a���p����^ ��4�JX�x�݇�Yk�p�˶�2�i��y���4� H�\#+�J�Ů7�L.����UY�:N���W:)�R��q'�z��܂���`�m�'n�`�EmMW]�C�2��X�=	�o0D<xo8?T����"4�s� VqT�v��#��YO:�o�TEE�̀P���^GzV�YP�COփ�N} �E�"]�)x�agl6��9o���W��ܑϯ$��O��8-���eT�� 5O���T�A�c9�q�,���r����*W�s��iRtZ���ռ��"���� ��D���+@d�gI�|_ѐ,?����g�(���X���=��$\�}�h�N�͠��CˇBe{��!�����T�n�Y�p�4B��d�E�kF�ݐ��m"�8����U)�.�G��B}G�g�Y
qU��F�F;��L�rK���B�M���Y�!��J�h�2�-Iƒ.�x�ϩ�%<��]�	<!EI�%�l$���8��%n��u�P�5��Q����H�+�1��;�H7�}�E����v�^��\��~���R:$a�b���r����_��T��U�)��4�G�X�N!v:C���I�.U��<���HE��~��c׉�-��O;�V�#�A��Eg��	�����`A�V
��x����j��P�9c�_��ĠDk���z7%M�OE��۪�|rd��5,ut/�9X�Bh�^O���]��������=���Oɠhw�A�������`'�Ի_�Mٗc@�Wto��y��X媻�
m�ki�9���g�nRe"�l�!U�6�EFs��G���^�8�dm6zY�-���v�����Q9@;ڒ�)M�^���/Tf�o@��;]x�R��J᱖|��l�ء{I2�BDXB��@c �
@�q���;��Lh���:j7��{��:�ߐ��8�����A}��k�b*��0�Yq�Ҷ&B�0�q���!ȣ��$���� fG��)>����?]1��z+���ǻ�nB~B<
��C~?dB����֮�j�l"�;���;�h�a.����������}u�A�u��8��|�.�����[
��W�J�~���ud:;��3�<�R���Ŗ���ۣ�N]v�1�?0���N���2-��� h]�������:�X/�S_�|v��p��xL�`�3��C�>ğ	f~6i��IL�ƍB{ϝ���VK���"[ �U:�R~�=H���*�2�GQ�ĲЪ����LE�V�3���;�쳛0�⼇��-[���g/��m�"�a��/7�-(��v�A�-��ʚ*a��%���IH���wPШLPŒ.�&��ߍ� ��@���/_��e���Q���P��4�$�&�`;`L�Q7�"G�H���R��_UCt�v�"O���Y���u/�;�wk���3(�_�Kq �}��b�_W���ņ�@lJ�.!�d����*\��U/ X��'Q.0�L�]�${�r��M.��:����wx� _å�V"Y�Q���G�,KN�O��Ca�V��`;N�g�z=+tJ�-�2�mZ�Ac��Z��\͟��ѓ�N����� =PkF,U���(N��5d�:ji�Ui���k{Bޘ�i��yC�3�[��7e�����0���"
��(i�v�βK�`/�n]�>���{/A��G��5+�����1����Bo���W�?�0�G�Pd�k5��)%̒1z i:	�$�IKFSͭ:nl@��o��^�B��: �~;�@�J��t���_�K����N�g���&vH%�h��'�?~�����0z(�#�҇�b��J5yXiN]��hW�u��F�6B9g[��5Ѹ�	
�}T����x�0~�m-3b�[��p��Q����5l0���9w�߫V7jՖ�o��c:6BA��*���6�q�6�^�1��֊�onw������"xpt^�Lܰ"p���1�c!�7%��{4�E9�*z퉘_�T}R�W֌sG�I_�;jC��U�>��>>5z�V�:�,Z���w����y���h&��,iR�����j
\��c�)Q-ݠu��d��w���x�v,�w��B��N g�n�3�2�:o!S�QɼU�72�&wQ�%� ,��(h��#R��0o#C��)sý6��b�ⱜj�'߁���5?��;����_H:}�����������y);��w�N#i��M7���z,i�?�T�ȳ�5�ud��%����^��,����O検�i��X�̊�"�lok��:/�-Z��A�8Ysi<��x�NҒi7N���A\�V�+,���\3��UYR���A�<KN��bx��������D��2L'W9�p�ő���
.��~���Ƿ= �(oPn�Q��S�u���aX_}�0W6{�-����H�IN|��HM����1�R)����Hk:��Hk"�3 ��*�]#U�o�.��7�m/ �v�X�r r��� j���.�Y��N \}Bl��[0�Z85��r�Ϊ���t�=��3�|A,4�+���~�_'y�?W=���+W$8C��b�2����J�s�zXd����ȿ���?��� ���ζ�F��xV�a�h@ut���ǘC�ۭ��!�U��qb1<T}��.&��<��3�zq^?<@��������YRM�֑�W��*^������?HϚ��]��%Ӝ�I[�����Mz���'�R�����RCWM@�@F�'��ꨱ��%�X�9�G��N.6[\��0F���}0�Ey�=���/_Rb�߅Hz�|]dm�lkk+t�j��R����Ȟ�Ӎoプ0��w� 1������1����r@�SbF�z�`"�R�Q��{	������)^�Y/��:;>П�.
�D[���h�v�3�����]y(ftr�h[��4G�Y��2u��e���P-
+,B����;}^�x)v�o5{���[iyY3�ދ����_i����6����s����U��ƒG�.Ԯ;S6Qh�%I�$Z������(>�<�H�6D��	�Ñ��7���t�G�[����ZNd$1�cJ�=jv��;�:}�w�G�U�cap{��gE,�5�v.j�d��UF/<�!����F�ْd�6[J}�Y��dsp��_����Au'��J1d�*-rz�7�W��!�U$�oW|�~DM[�-�a�CwJO���w���\��
��o� �,GP�=��)��_ȣ����Q<��p�v��h���~�i%m*$㜩>�\��
�o�)�PP�`����B<z��gT{�z	 ����aW�G��4M<������$|�)�W-�-�C�¡|�%�.��DQ2���N0��T>�A�'�7<=9�L	L��X~�rΑ�5*����7l{��U�&�O�\�m�����^61�qm�Χl���ͮ����~;69jp�V$�]�>�#�� BLK	Uヺ�\���*����@O��p�)��r����44H�Q.��2c��@���E��5Hw�X��^ghF"���s��к�x=
���t�\Y\�@�w��0����36�J$��/Ѷ �V�;�o�sAN�R�S܄6�45Sg8��T�0��v!�bl8GH&I�e�dj�%AΧ�и��g�)� �3�����->�x�(	;I�qYܰ�Q�[7_U�������CR��4�MD/�'Y�ɼ�t��R���?	��Q�4V��	����E�����F��v��z���rY��Q/A(�W���<΄6��u"db[̄&�ۯdl��Y�FOm
�
���Q2��[�K�l a�%!�P�[�Je����s�1���������s��9�z�;�ͣ����;��B#���3�2?�g���wMy���=��a�ؽ��i�v|ɗ��08��:�)�t����q��b(~uo˜��<m�36�bU����Z?�P��J@���O��0п�ўqԠ���!~n���#H s�f+��.����^u��n �v^˶>
R_^�(��`T���Pn�d��ɩ/���~�ȫ����YHrFzG&�?J=���.JP+I�����35��jI�Q�Y��l��93��@�L{׽	4�X�ŋ�,�{��P�\�'�+ǚ��G�7x�]И3qJ�c������(f_[�`�����tC���A�:A�삗�<<�a1��O�.���-���cs�5P��� ��	"�d�nsD4���6D�)�������@>��=��y�2����I�O��Cn�j�xP���p�8���1��N�ܻ��P������x/n�3#н���4T��rr鈍���ʮ�xж��Q ��	�_�#�i+���i}������	o�>���#Yq��>cTo/g4��:$��n �*<���Gaߞߥ�Y���c������ly8�XVO�TN��[a	տv������6�
[<�A ��6�fJ��^�"B����h\��M�J��1ί�!�^�C�5�Qa8DIlND74�����a)+nl�e{��%H�Р}tq�=���
�����T_ H��fGBal��U&�8w|X��D5�8	��a|�Ay���� ���)���:�����|:�����-^��ڿ��,�S�� ��f�
�Z��ɘ �ÿ&�Ȝ{Q�G׾�)���8/��J��.�+mm��� ������W��3�J���S�A�] (���ń��Tt�)�+��.�������^�9�1�J��ʵ�V�pJ�=�eu�?�t�]�%*�O����:�Yw���r�3I�=���%�yTM.�M��MR��2(LAg��~����N_�88[�53��T�¨e���I��n�����+�0-�b�3Y�\lGn�zRY~��Q2��d�*v���*�w�� �sC�.<�O��������jyd=��D�[+&���+#�km"1U�&�����~��66a('�C�Z%}Ȼ"5抡������52 �!:gƹ��U��(e�J�qJ�7v�+X�$"#�|n������ζ_�E�/e��ȝ6?��IPR��cؖ��lQA����Ֆ�\ꆘ��������w�A�S�KO`S*5�$�ڟi�;~ת�x$1��"�0d��G ��K�.�������5�`I��*R4Em�������u:`�G�
���o������g���J+EqF9Oqw*[8��t���O�y_RZ'�.Fc�r�ldLu���+�Kuj� �U�}�ӡ�Z�
)y����RHj�-r��p�nf��*�<�aQd���CNL	\�����  �:�Gq�f��" ��ң�sq���${���w�K4���(D�-N���6jv�����*8�ěj�'iC�����z��5�2~��p�c�U���
6Fd��Y!R��c�%�*���fR�d1"����%�/����S��C���)��-x��@N:�V\��G$�:[P/>2d�ЇVK�U���j�"�!5J!A�`-��죐�h��>ZƋ\�zC���1s��M�8�0Lh�`�o&��Z��ϩ�E"K� g%6Q	b�O���_�� 1�J]4A'�%d�J�T���U|Gl�! �w��p�RB��%gf��)�b�SLv�����
Wkc���>�c��t�>
�i�J�#�7��C�oD��ΰ�8� ��)�U�1�J�Y��(�ez��6���:�j��tL`�u����i�=Nq���TP_>x٦�v�$��Ga=�'�:Dc��q���8X��P�Ū5��>'�Kz�%˲�=�V��8(	�����P��D��M�Xй P�I&B�ӑ\>�g�2�]m0�>}���D��y�)E���.�B���6]��kV	^m��v�Η�C{��
���1[:��BD�I���W�ڀ�	�_(�(�M(U�i��)]p����J��5a��V���t�	R�J=l��H>�:!d����-���t�`�����r�e���zQ0H��D֫�N�g���T&����\�r.�g$�)�