��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���!<So���2��E�!�7���feI�R�34�F�\1uR�XO.P㤳��"����(W�����Y�us�'�V6g{���/�Y�^( ���Ne�[�����8�1��{SZ�k�eZɇ�FUHn�i!�ӣ���)K2�`��}���Z��ÏR��Ȩ��՛�,`� >d��XV�i��[�ss-���\�Ж?��麱t�/�:��+yaxp;r�V�}�S
ꜘ1��y�ar�}ٸ$�	�"�P��Κ�y�t�s8l ���DV����Wi*���
�> �=�IdG ��Mπ��O_�v�����?�m9�b�d����k�v䥹��/��֯]�G�W5b˓�G"_?�T3r|M�u���j��$� �V�p����"4nQM��Z��7�n��H�E�.G�	MB6��W`�>A�k.�G������q�$p{6�b�U�Ϸ���E��D�P��zb
���5��҇@����9���'QU�s�?������[� u)��4ȡ��S[���TpY-Bk6T�B��e��CsY��)%F��/Ķ��l��"�WA6���r�-���RC��\����b��M�߇��%|�ɗ��n�1O�f4q��=�7����":x;������,Yv����{��F:�2�4�B�N��,=1�@�Z��Cōa�(n̹��Q�ttQQ�_X���H�`8���2QjyT��[��E�l��ʌ=���*L�y�NP͖�t�3��E�� f�KH�Ɂ�Z��g�������-�&�Ȓ�Ҥ�H��;)�\�M�/".�S=�r�鱔f��E;
EHY;?{�
 ��K!��+����sm�e �$�/a�>�ى��i��xg��X�'H�eW�>����![y����0r�
�Ac�R�b �K�]	���T���^�s������'����<ؕ�w�:����N�	�W�p�g�*K���(�6a����cXa�.J���]�1���g�]�l�u|ֽc�)a@���Ȥr)���<��f��������N���5�Z&@�l5cR/�ݗ�0�����>!�	�r*�r��aѸ
_2�| !�>����M�#$-C�F(�� 	/���<W)�Myh�����Ƽ%��E���j��>���nܧ!C�*�vkH�d�(��u�J��@��F}up�*K����W������o<]CAMw��ӣ��衟�2����źG�.	��C�h/(���������^��@~af�iq�L6�^0�Շ�׻�c�~�3�۳���W���43����" �c+��b3�(���"����ix�
6v��p{D��a�a5Qn$�S'Na3�K9�B�b��^g�0���Y�8���x�q���޷�YK���L�q�֡�	�믢��r���O螊����wN(9K���Φ8~_�/y�S��>A{us�|{c��3�8��
׈캗�ڒsn4�I�)���r;���<�_h;��47����f�m�qXv��o<���]�8�I🣋ڏ�03O�]��Z;8�?�ŢL��t�o�nQq6�r7źI��Gɮ�a�N@{.DȻ��͸�_�����3�/���9� C����,QA�,:�r��ZQ�J:�^��k�/ C����C~��N�೭H��H%�Z�?Ɯ�\'���tI=��X)�u'v���:���l]�s��v���}ڟ1`��iʂ��+�&O'��d2~�`+���̫M��ek�M��,q������M�S�-���ѳVc�kOc��U	����2�_�A���Ơ�E�����ܯ0�< � ����C�Aɡe�1�n#Q�Mّ/:(���S\�8��
�9K��k�y���+�xu�\�]�m�����iX^�f8�l�#LYan�Qf%-�n���r�zs֧]���D��h:��{iR��v�z�)�;���bDI
��ZKH-nu��U����kf�,�FFh$4T
`;�|.�������xm��������&��T2��V���HP�quh�S�A����X(�n/�%r��/,��w��!%�,6������׀$�B���&x��H"��E�vZ00c��;�6�8_!�Qx]�a� ���	/�Zn㲄ôw�L���HaN�B̵mMk�d[��B��[�,	�4 *���6���ǳ,�҉c>���]���\�;�E^'˳�H�g"���r;�]��"�t���E436�V_�7eh�4

�qHe���7*�۞@x ���}"�#�H�����l�m�#���+�#]�ÒsH���gî��|�>=l؋�rb�CM+�~CT�*�;U�'@e�H=!2��W	&z)�t��*�����2:
�d,��ށ1��`�'dRqM��,X�f�;���KR�Ԙ$�Q�t�>��鰴������M�X:��l�H�/#r¡�Ԗl�N�"(�m�Z��*��Qyk٘C��<�C�Fo���(�sJ,�oh���~Z�x)��T8m4G3�ct���Y����&���~o0:kҐzd��A2� ������h�U�s@�<纀pm\��>Ԏ�$*�#.��c��Ɣr�~��4G����2��,n�|@l����XЍuѾ����H����u����sn~��G��Q�l��[���P@�,%��&;��"�;�`�Cףru"�Q<oL}�ٶ�'�9�7��Kp�A��e؏�z�ԭ`����Y���l�o����Hu��A��K�{�0�Z�&�fS��L,��>k��.l��%���!1]�{���I4�Q9T(HSǫ|��1u��s���S��s��e9��p�@t�ƉI׏�Zֈ'�i�ѿy[vh����K%������-�"x2����F"^���}gg���IN8c5b�lpH<���y����0RWLi�?�w�{v$ܽSkC�ڡGfb3��.�B?1i�m�f���}V�x�W�=�VE
�l��/��p�wĘG�,�9)}�K'#ra�����f��-�68��I��U4��=g�@�G-(�itz�ҹHt.�X�:�4r�{P^��4'���~��+��P�2W1=��t�\�ͨ���k[��H��G�,�QJ�Pc)Z�Ȭ�'Bv��U��,$!�H��\�o"+JN�_Ҫ�=�&��>���-G��R&�6���_%V�+s7�_��7,,��6��i���}`�j�2�9�x�` VCQ����������ߏ��;�fD�(�,����������W@�J ҟ!�H���S��f���A� �r:oh��6���6�G%�9��c�M����^&=�^��7#0(���߳]�����MW%5��P�&��6�r�|��X)�0yC�*y��5k�-<;xi?�����CI@D�9#��N;�:����i�|_�cV�g������$���e���S��6P��o�0?�����	�����m�/K��[q:���r�cm�g��#OW)�:'Hވ�L/BL�#0�IV�>>`TtLq�)����G�j��ΩV��fq8@���X�]p�8!�D���B�g7%���{�ۘ�F!�ed�{��ߨ�2���ô�S���fOl����7�����:�|�ʍpf�@��o�+���d"8�2�_S��n-P3�Y.��i��Ӡ
L�~U��g��>}����3�Yވ+�#���Z�o�0��0������N��I�V���G*B�>^��c��w�����y��'�I�X�! B@�E�p�*�.n�rd7�oeͦ���y�����<d]s���m6���y��.��1��0��>��z���S{�G���4���/`��!u�+Q���8�A�7x�Y�'RO.-���`�t�P��2җ�J�f����x�BTE�d����i�D����}ۋًsT�i;Ɛd�S�R9���� ��Ƴ���l��[�Q�c�d�9������o��ҊH��O"H6�Ob>&1޾Q�s�-L����I#$�K������X12�Lq
���MwA��hM��?r����<�h���c (w����CF�4�K��<R���(=�J:�u�8�C����T�MWiV�-ȳ�$��Wl@8������u��F������#6�����D�Sbz�JT����������z��Q�V���	��y|s��4�P�`S�oEIN�kk����+��ڲ7�i��;��l�`Pў������
k�UP�
�o�;�Hk*�4S������#��^&G�;��3��"�簛2l��ktJ�PBАJm���1������:�{C�b�}m��ߑ+ՙ���f�����Ɂ]4�h��J0b� y�#��sAȕ�jLӣf�%�� @����w���4)�o�zD��KZ�6�)S�0��q^:ik���9���$'���B|d-SY���鎁�t�G����'"CW7F��FZW���J�荎9��֏?�u�R���|�8[���A*�:����J72��3��ZX���^l5I�;���s���y_5���R�O�������ح���=�4�R�x��ݗH���zY��`>�Q d��&	X,�����{(!?��ޮ���qޞ��w<� b����+3m�@���`�&���ao^�����n�Λ����*"����xnTJ�m��I�(Eڸ�@�}��0�xmar��sh?a��$��^$f�u�>�� eԔc!6���y��k�d� ElZ0V�D�'��0�����Y��d��(k�ͩ��77�����{7f�&1+���G��]���g���P*l�l,�����^�9�4D���R���v�Z9)�O�ױ'7�5�Ϣ-I�t��<�&���:7�8��વ#�ng/�uS�Nræw��Bp����u����?������$��gp1��L�AH�u���~N�:��a��v����1	���������Ť��7S82��+���h���2�wbVX:�r��x�=�@��n��,��}q�L����z����/�P����?o]�H��6܁;\2V��yB>ak}L�M�Ӟ�N��������b�a(E0Iǎ��kN���g�U�`�،np��;�<V��v��G��Lݜ@{UJ�U����8�J+��իv�}Ҹ6���Z9�G�aN�3��t�%���>x}y�����Q(8�~<>�l���%����8��Y(:2�J6�Z�G�o�WW���a^J&���ݢ�o#�ƿ�?��/y,v��}��g�C����P�^*��.X.��0�]�ڮm߸�K,�Q�d�:곗�'�j��`����l�i���vZ|��� e��}!�>����,��wb'�)��n���g����g
���k�����2�um*��j����>�tC Ͼ}!αr49��c7j�|��~��}��ֲ�~�"Ԑ'�dϰ8�:i�ZiQ�$�H�(Ľ�, �8H�.��2��h����̓}��B�!��2�}��*^�~��i�1L�B���e����J�<#�3åv?�=�~�9�^�*fq"�+������ns�������_?�d��e�JMN=�����񾯒;���Z�i9���ڻ})ux��Ϲ��R7�sE�%����u(ud���_��CΧ�ZQ1����iz������Y��&���@�/nc�F����Gb�0���$�}O�4Pp�j�Bt��T÷���o@`�R�['�dR�h�)F���2��rf�����`Z���= zb�!T�l�v"Z�)�jgO'��]XRq�7�ۆV9{ϟҒ�|a�%�.�t_��+�w_�9!� �68�*�G����-��e��̮@[ ��z��!JI����{��ﹱ�]��/��
?4#0����9�09��$��C� fAnO�K���{�����I�����|�v�dvx~(�E����#�WV�����r#8 .u*[6݊g�s����~�A8Rރ� ��2��f�w�����yR��Ra˩�L�؉�������!���Z�7Bv���Q�)�0�)OxT��W�.�GB	�S�r-����X �݌�������4-��fV���$4їtl�P����)��fB:�s+�;͘����(��W��:Z�P �"8�D�2�����K 
!+�L�q�/2p˚u�T2�w&���N$A �>����}��/%���$�����*"�Y�{̟߇�i�J�[ L�'��D��b�o�t0y��	SY�8`������g�k	�ӄ�dw���F��(bS$�� v�/�1a�\����J	��	��/�T\��a,2�,C��3^���nH��Ul�;�Q܌��mv��C$�>V߳ԍ��"��R4J�'T���k��a�8��W8�H�.�K-� �x���x0�������G���N���H���1].�#fl9������i>��N�\�CwfͶã���^�*�֜�u4�<>�T�H�<2�����V�O�a���~��g�����p~xԁ�v��'��E�#!�A���	B��� ��)�3�-�4wU-�?D����G�[ِ�z
�`-���]rz�>����(8`�Ζ�o����;��u1�6rW�E�Ɖ���v���3�i�qy������b�E��p�o</ 9��y�����/�\�r'�N/#��~�t�F����B;m�PW��,�ҳ=DB�g%��=u�M��Q�׊�-U�>�̏�*�DAn ߓ�Gǉ(�"���q�Pܒ�y[�Z��mX��D^\�����������u0�'�g{G;����;�h l*��~j5�\�U4�~S���������2��M�V���q���o��B����˸%��z�k��+�����Pg�Ĥ+�4ec��S.~V��-=�1��U4!ޗ�L�[ `7rUjph�^�k�	"�WY�)!7�oCd�2KP	Nԗ��~^LQ�������\�~�Ls�%7[N��/G�s��-
�P��Ks�;�ն�R"
ɧ�W��#nߕ+^�?+p����hA��?�v�ڊA�|O.����t�f���@��_Y��/it���D�MF^!��k
k���-��[L��R�������7^p�Q�G��M��Ŵ]PƩ>q�ۖӺż}�.ݬ��V@n_�	Kp:���xj���pO,X4�;�0N�^i咼a@�lL��T��b@��̇��q�,5o�┧�vyZ���ɶ�v��"���e�S�]���ԷmYn`9'�V��Z�Y�Z�:��|W/i6/��$���3��P�zY
�*��"7KAH?IF�l�SS���I�"��aem|�B��[j�2�EA��#b��8�������D�, ����V.A�8I�8�M���҆]�b`W��`s�x����*�ڻ�9B� �>���'^�#`�NecWֽ?H/�Es��5}�����<����	��V5��?6�sɕ��6e�)<�+��-�P���Ao����ֹ�e��B���l��IӃ���)��uW�9��e�J[��š��8/"�@X����PxvyEיP>@3=$#3v�jw�������DtH`>l���w�$��y)��;�WuojlP`�Fb�}ā�c`�Siulb�
�z.��&³��~ n�N���W�8I1g��"Ri��\�"b0N��ȩ`VtLӾ�K�������tt������F����Ӈ8~�y+��V�Y���>��@��\���^�]�'�lZ�A���*m%�pu��)w��\���e�,J��K��g�A�h_#�C3���c6��#N�>����3�˟�\��[a��b"���,G�&qT�GU�����Ɵ�@N��(��)W��1x�p��3��-�p=�SsV��P��K*����?����F	���*U��j�k���&�f�p������RN�[��5�u$�����t��B� MR|��@�Ⱦ�6Z���:���+׎�R�DlѸ����C�I��n��>ؓ��/������P����#����J���f���F����?�ö��;.P���Z�eu����e��N�TO\���:��4oP>^k����Wv\m�,Fw��HE��12TH�ŕ4�ikO�p�I�������/�	sv#�t��T12]~ZH��I��3�gu���3��P��a���pEt-���,w�+��q*��ڬ�L*[6��zt���Vÿ�``�}��9�T%2���i�[y�!�!��q�v�f�<��,��ـ�m@mi}��c=��˻EF�O�>���x�K���c����y���U�Ұ'\����� �$�g�5�Y$߼!�ܷ�� �M�Y*b;���-�V�����Q4�Ż.��{ѕ� ��@��l�.l��/���X(/D��"��`��H(�׎�sƢ��͉xE.X�_WM�ZSo>r�,�e~�%�1p��������T�)]�D�;߮�	T� ���R;h$�Q�`�H�Y=@��2�o�+�H����bRɍ���$��G5�W�`bזn�f�^.���)_�������f����ܪ�̃����Ö����O�L:<��9ghr�B��R��V�,��Vt��!wh� :sNS��P�M��:w�����jq���U2�WJqMVa�N���9b��̬O<6m�*�!Xd����g١< R d�@>���M3qRy߭^��Ǌ3�|�b~M�vZY�_��ԇ9������'�=��d ��f\0�{~�E:5֟�F2���gMH�O_
�!���J�T��x�cf#"Kӂ�L�'����Kֺgw5�\����]�~��W�݌uE�E>�LD�
�%���l�t@TV��PCLّ�;&Y����ӧG��/
 =��м��[衔� ����y9=~�N�����͌�Wx7���T����g� �Z:W�i��\�����?C����R�w*К�}���^�΃��h�8���?�b���Gb9��z�j��A���
�!���C����(ХnZr�bR�.��Ǽ���:�C���u���av{s�DiW`V��`����Q����T>��B�	vaC|�'�2�L��t8l�����_eAi@��!�m���K��3,:�-F���Տ��ƕ�����B���SvK��/�JG�����	L�;j��'B�~��!74�xG^��s�Q�"��,V2Q�ʇ��~>}����.��sJ��a!䵯��^�K�`�bD޴N�GS��on�i���� �&`5��T�y��b���wYQg�p� W��С�AJ�Ţ�_Tm�R'(#�y=C��J�����v�gc%n,'q$7
/w�V��QR� J54	'�}c�%$�{Pi졻.}AԲw�0����U�biG@�n"h��Jj�!�y�a���W��*?	hs��JfuZb��Ǿ��2�l@�_u���PM�qQ��7p8����#d%��yĤ8u�'G\&��Z[��~�n.b�.���Z1�!�O
����%ڏ|�� ���"%�ӗt��bR�'�!(g#��H�վ۲�@�1D,�v�y�4y,��g.4�����\a��nM�������0�߬�V_0UqR��ū�I��4�h-�:��'\b���̴<հP��6G��1*p���\���Ւ\qo��s�j�#��Y34��]5�Y����:ˠ�����5��%����m������0UpLFtGcTy�P�@/����i�Y����q^A$m|�~��i�)-W��f��[7G>MQ��w �'�1���ҳ��?�L����GT{C�%ҷ#����^S-[�����<�ĕ!�x�s�4�Э�]}���^�F��������Lı;*o�.�_�'�j<�\\��0
_�N��ּqe�JZ���aL
h�rl/��e�{"s�J�����h��$������ŒMJ��(��>`���0��n*�ŀn"É?���?��1Q=@�h���Ts{'5�x��4I�t�C����+r>b�
$s�}X<�,!8����30�=O�������{��J颗b^�{7�"W�Va5�����T�����>ꡭ�q}��G�W�1�&{��t&��{�K�L��� �)\)�uJ�=������'����7�Q�YQL��`M�EW�,ٯ8/8�h��T��?j7��/�����<��Cp����!y �XWV��R4��ļ�OuG%{��YCY�(+�q@"�K�6�)�+�3�5����N� ���关E�W~��UeF����� �q�/a��'��s�{uȾ����^�l��4��٫�}���ӡ%�w�,��
��x|��Y{;�;����}�y�\�҆ϲ��Q��f�d5Y�;�'	�״�x�]�,�:�D*r=���ڎe&B�r�# Z��Le�>Z��!ҠD�S���#`�-�/�>�Y�i�
��?��0��		e�Eꇌ��Cn�o��GB/7G@N"��*��q��R(!�@±�xO�,�ѕ%���u����/�[�~�p�|��~�Ë�����|UU��g��ަ�1�*|���<+^dĭ�{�~}�EG�V`I')�"�\�J3D�IU�s$2�%2@k-@�׸�R�YPT���k!�����Yr�����lAM�T/���C�knJ%�.�7{#�}@l#�/��~�}#F
�����_o7�a�	��l&�����)�	.8�E�{�ô����u�
)��ؘg�U�J$�],��|�mc��>g���*!���L����V���L��,��R��o�P������t�{���B���2�u����d����<��o��c��o�y�V-�G��Ao��9������1u㋲o�kHB�2HPo%���溯��P�Go��`�����L֏�ж�c)�S2'��tW�t�Ȭ��c��2��k�ib{d�G�1��x������
��-�µ);�O���SB�%|[��t�bL���\����`�6Mp��LTȬ1C����Q����2��d'��S�,&1�߸���q%~=��m���Z۳KP�1���V2�>���MxB��Ȥ ��F.������6�?�y�<�u�z8bS=����U�m��T�Sj�4����!������󅯓O�A\���E���9P ����/H�`!��/D����{�К��v�H�vo�CVO9�kr7`������(���_l�3�g�hr�jߞɘ'.|y$Slί7��%�Ԍ����?ڲ0w��pO]Bz��]d�zWT����;9��`���.mh�{q�8�faDslטT�����-��gl$�J_�|d�+~ga��Ӑ�B6Ɵ����c��/����*'w��Κ�?d�=-v�l��51.��YI�ߣ��¬t���:!X$�7X5��]P���P}���ܬՄ��+GC5g�z�2WTT�q@#\������a�W�Dx�i`�/o��0	uϝZI��I�L$<ɇWZ���4��r>\���� @�|���e�T��:��bO�`ىi̯h4DI��o�s��R]6����
�bi��z��I��\>������4w+�ܻ��W��_����A�`���Z�B��U���v*pH7$�E��4��攞�kt��%�s�K��ߥ2��t3��Y���_��oc�[��D&�0�W�H��?o�NSl�O�T��2���AL\/���j�-���i� �ɷ�32�M
���yQ�G>@\�S>�������y�������sn�݃��X�W��6G��xҌ_O�}:0�{�"	 �_s%X��?�����W�,D;&8�y�Z��7�
'��ħ����v«����^.�����#~��!�3A�W�[����4�7�� ΩDD�Yy2Fs��{v�u�i6zs��r�'�����)��
�JdJ:D-TR�a��E��R���޿K[.O�L����[��k�+�/=�> lI��Q��F���(�{x^܁�Y��Ƃڙ�N�U�;.{��3��'F������*a/~���{�C��5z�g�M��C�]�d�q�o��ȳ�E,�s��s,��?|�4��*((�
��'�vQ��}�b���tZ�H|N0�am5����ҩ�<�"���w��s;;#��~��vo�h���&'�w���w�XLiu3��z�п����<�O�q8� �-$E�9��m�<N�b�<�
J251"&���Q�gÍ[?Z��Y���N��޽�P5�oJ$k-���q��.R������3U�/l���6��ES������+�9��'�ս���>�/�i������Դ�c:Em���L ���h���S9���9xg������e�y&F@�u��=�7��̈���M��J�+�E� l��F�m����b�k�F7UE�U�/�N >�sUvN&1��:�����m�Bޣ�Z"�� �4fV�6�u<@�~Y�8�><��)ս�I?R�un�x�Kt���2���e��*�JT��&��7Ң��Ҥ�߼��lۭ?;����ә�^V���N%���ШC'�)���Y�� ��ٲ��s�U͖��aA�h#H[��4z��|Dc��T�f��b��2Y����"�G��jH%>U���ѣF��0_��k �[ߵ��F�2!/��NQt��Pgn��w+vY���9f��þ��/�2o#ɑЍo"Por.Y:���(�M��xA�^�=Q�ģӥ)yMX_����叶%�ӯ�ʹ$�Ov5��A3��+�&1V���"o_�����
V���u h�}�t�9�{%����Z�z@̶?�����a(����m�b5z�J�����/!���)ϡ��	6��ߒ���-j$���=0���o[փ�!I���XE��duV�I�߲/ȼ��w\�e��ﮆ�k����6��ҋ�����UY�m���k�i*�w��gR�¸?��y6�mG����،o�	�����_Ә�#�O�1b!�B<:;�MlV�qbZ��A]O3��1�����qZH��3�#�����Z�um���s�t!�@A������O�0�שJ�)T�����3��bؒ`	����d11q����*<F	`Q#�n'����Kޒ?s�T�8bT*����[M�%�W�T�@�
_���ɔ