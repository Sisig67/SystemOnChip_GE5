��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_��՛	�D
������Jl]Ǵ�j��MioL��
�vf���~1E#!�6�_.���㋟#�T�Aw鲄���*_ kf�t�:3�٬��S��<�4�O��K��v3��_h�W$*���q�7g<W����W��ԁ" �}�%��/ʨ�x�2�HY�] gS	l�o6�y<a��Y��u4���x�*JaSL��&		�Qv����(�&3���WZL��B� �)|�T�����6x�ǰނm�i��Hv���層�Ǆ\�On�= s4g�J��<VP*@��uκE� �A��h��*6����Qm^i�W��5k�[��:X��/T����h�j��HP�ޑ#���.ؽ'}dodr�qK-1"_8g]�6]2��1'�����M�0�	^_�s#�j
�<�g��$��;X�g�B1+���t����d(3�Z���ȓ��/��%��v��;�Mo�M�h��?���,�B?��- ���8�?e�V��d��E24��������pBz�od0�q=Uhu�����*qw�FcmX�Xk7�m�g�Y�1���%�{m&�#E�kq��9�
�*l�!f����SP��)/��&ꩥ�����L2KMJ#�<�I}�D� ���2t1�C�hU,k ����l`���h�����^>:�pK�]W�\ű�[�'��V�O��4㶇�5��]L� �<Q�u�:*�t�����!:�M�L7�!�R6�r6u���D� ,� ��s,�6xߪ��AEt���	�>X8�$�������fdTP�� ��L�h�.�o�������6���r���3|��Ba/;�s�ڤ�.\����e�ZO"��j{�|g�M.����g��p���.V�2�-�G^�]x6>,� p�  6�f�z:;�%�=��b��Ì巡�faBX���z&����Hu� .��ә#t:^�ӟt�v�fG}���n� �g{�LA��p�g��&kK ���Zy��Tn�U�m�'���
L������F5
#���U�ﯲ���M-m������[J�lƞH���=�\ҷH�:2Q�.�<A_���+WB�� �p���9+����$H9��z�7~
�+`w���	�5t�KE2v#f�d��C�^3/�]%нP(),�v�v��^��װ�y�s��;�E�SאZ�U�хf��I����+V&67Q��"�
\uq|:eQƺ	8��}�+br�ń>��& �M��[����m�2��2�L��;$)K>9���P��Z���P�����W�@��G�ޑ�7l�\a�n��`�"R��,ŭ8>����-�.#����B=[�]X�,�\�Η��S�]�ҟ%���n�������I���Lդ�Q��(N
_ �3�Hճŵ�z���g���8��K�����!�~�X���O��s"Xw_�9G#���	o�PQ/�K�#T�c�뿜��a73���v#-ً��Z�zg�|�}�\J��ӟڔ�\��{ot���G/�
����ٌ�����G0c��	8(���e�|�Z'���l=�b��p�6�_�7xB5��`��q�p3�-pD��B�|�>�\	��T�Ѩ=����`U��>��&��Oc�v���ʯ�8b��:�<NR���(�cOt9��#�,3i`Ug\�CjΞ�!������Xz�E)����K��^:��.�Yit\��<��1��D���{N���
�׍��.S�K����oD�K f�R�딬Ȱ���x��qh�m8x�_�g��'�0�>����h�����,�5a�B�ԡ{c�J\��K�S�d��US��i��7�($&KDdyh�	������#f�$.��kN.XɃ�I��΁�� ���>|J�n3i�pT[�O��r�?�o����8`�ǲ����6G�n�8��{{RϞ�5��YB��v�ReHMS<�3�b��$W l�믘��u����Џ��(q�I�Wq�'���ٍI�������Z��hܔ�`>do�ﰿ�Sk=�����N��a��u��P��X8�y�|���(��v���Q��^we�*��� ��f��F�1�;�JC�r��m)<J��j��Fqʊ��h��,4~'G�����A�[�&��K��x��<�� �` ��9|��)������P��%���N��r+o>j��X�͊ j��Y)\�G@.�Wy�[p��nR��!�F�0j�80N�g/�	�u���֬K������Uʕ%�]�݀��0���/�3��M!�%K��s pe�,y*�� 􅧶O3���I�D�w �:A�¢ �#�����i3��n32�5����M�z~�ʅY��8�q�K=�|	E�RkO2�MK �V�Q����3sv�W� <6�z�)-\Tgl�HSD�k�~�\v;�_��Q@zb��*dC�ͣ�I�U��VFQ@�֬l�y��q�� g���*��\ۡлs�"��,;��+�	i��:s�d��h	����Տc�O&[�N:a�-�z'�_�}� �� u��0�v8�������U��/㲪����3�2d��)ΐ��)��k>��ٳ�*$�����$[7��[��j�=��M�o|��O���)��K<�/���)�'�Y2d(���x�D,֮{�i���'@�z2�T2�rG�n	��Νw�	jQtrE��H� ��-�ȃ����-[��iL{Q$)�j;�A����2��0��Mp��=�a�ޟ�Up�y3:��o����r������eW��]������&��e�5�4"�O��2����a\�ȸ���#�I���86)���O�X���3����'����\���U8����0>8Zl�Ɯ6�4�[Ӱ���jz�̀8��[��Ys�Oh��N���!WQZ�Qr�����FN%x��nM�ο��As��
q~'D�'�Z����������1��䫦}f͎���YC2�!8D�*���Xnk�\LL�' '7��tv�6`(�azT��J���FN�4����5�.\U5��H�	�LO{ٳ�Q!�3��~X1�Q�*�쏫�&}?����)
j���0ȯy����}Ϡf����@�kUL��My!��Hu�+�U���;1B:���z��Q���>E�>-��j��0�ݽ�QS�i�o]��>������[}��E 7�+S��E9��|,��n�iPZI����E�b��_(Դ0N�'��F�5�k �.)�\�/�B
Y<��ؠn�Q%赀z��{�M ���FV[P�3�J�X���~��*9��߰k�~�v*@��2��
�ݪ;�T��$��5�NG���Ҙrw��Y��Q� �5T=|ӛwʰ�9�u$��u�h��^��S!�-2ϓ����Т}^�N]�vC:��5���n �&;��E�`#���F����MY�|)NK��ȭ_�NO'������Z��$C��s�����*D<f�J�g��rCk��p�0u.a�͍we%"�l9�����K�,�NsdB��p��/��$��Z�Y�ů
(��~zo�	;�4�wc�,�F�?����(#���=�0���]��_o��ܺf=�Ž&9!]�1=U |�4]G#2��$��L��%�ꅘv:۠���&�� e`묊��1��n�H�nRG�P��z��jL�r��<X7��=�/	j��(���X���)4Rq8
݅�|�$^���1��3<ѳP��-�$>�*�NO��A��F���Am�P̘rK�U���3�<������=i��YAc�����id����l�2��qx��49�U���Lh������#!�F�+�A�e��]w�a-�W�ڌ��Aŉ�����!�j +�����yV��Oܣ�/P���4�8� �ZLP.�C�$����Ҟ=~f�AfeC������������t��[q�¨��D�t�64�����+253Fb��!��q?�� r`���'U�N>����"��T9%���F���5��Yk>1L.�"	7�xB\�(�-��g��h��l�J"��ٝ�R���8�0��Hxpڮb!z㧸�{�6����.�5��N_>��``Y%Ê9�0)��=օ� �bZ�M�� ��R�������d1�Rm�����-�ƾ��ԥF�![|H�o���d,��r�{�3�U"*�h>P$R��+qZ!���q�+XƆRK���/N���TEB����w�9trx��M8��܈kfS}��P}��oUK�K����Y�v�{FǵZnj߿U#u�o��^33��K$N��7ª�j��
�[l�q�gg�x��Z�|����*�Yl A�륯HOÞB�nz�I�~�@�F[����&x{��+u��E����i�B�'6O�: ��V�ڗB�`���h�.����{����(�k��~7j�'�6�@g�xp���:�2���AQ��{���K�;Z�⥲s'��hH����A��x��\��[��偏��(z�e����dz�e䅷ω"	<�d�&�[��^ѝƐ�X�?�>CL�J��d����? &e��:1۲A'Ձn�ѿaJ}����[�e�&���b��ʟ�żF����4���;���| j���e,
:J��G��nZ�F�B��
f���
�H���c:��}��\3.��y|�+�4��RޫʚQ�I���84,~��O�\Ҳ�9�B|��46P��Ax��1�M�/$�ʞD�Вy�!��j5�LLM3��G�R�&~��.��x�%�l2s���Ɗ(�@�v���#��)���1l».���)����oF
���n��' t��8��v(���Y R�"���&�
�8���3��U{4�HcG�W���O��R����e�����B�p�f3>^�Ny�_��W��P�@�j������+w3���z�>Db�h�v�(w��XDD>X!u��-��T�ɿ��8�%�,%D�����s%��"? ��f�i���	��_��9��CbeM���1<�伒�~�Y�i�T�%ߠ�`�f�`���*ʣ����K���^���bV����ї#��!�G��ɭ춀�������MG����F8�n�ݙ��?^A��cڹR(H�NBb��=gM��<l�K���!S���L�jʬ�	tBr�r�,����o:bF���W9C��	)C��*I�ɘ�S�yp��F��ֲ!�#oS����+$5��3$Tev.��C�[�?�Q��ܙK *h�5�NZ�B���`���`��ib�E�#��7��Vk�$������z���|�npCʣU&\��6lFf�=o��D�{;@	�1�������@=nm��66~VZ�n����դ��|I�I��jr(��|��/�.+��²D�[�:�;����� ]x���F�F.e��|k���@8������aXc&���!z�O3N���d���C"�T�|!ڝq�6sX�����.+�g���ea{�v@���sK��.���@C����Mk��'a��$0�&�n,3�v��Rc�v�Hv-Uv�F7��`�|qx$ tָ�X�	\��L��Lwl3BN9B{S��@�h  �ᾄ�g4�,|��L����FkN��ً�R.)�E�6@����30�����L��9�	?'�Y����Rl=;McXH3�)J&W��4򥥯oF>�q<�#�� p��bV�	˖q9���X-�0l��b�B����!3����rɀ����dnW�|��5D��FSٓ:�[��Qp�����8ҝ:��٧9��i���>IN(�Md�m��2�cvj73ԟ>([x(� ��E֡v��Q�he٠u�)��x��37y3yg��s�8JÕj���I��LE�\�8�@<i,p�W�Dp�����5vA�v;#�b��H�^����l�M��Qn���
vL\6;d�1��Ҿ��F1#I&/oB��u�2�uߑtn����R�83�Gd��~�����U���n�<6���o}�P�I��Gl��	��|7HI�{ꮅ ���A�\��VS�0s(�5���ZE�>k���Є�����U{���99�d�d��$b��]P:h�G'�	5F3̢o]WMy���*�s,�	AG�����GԖ���r��F6�&���2�UEB�f�
%qE��b@KЗ�6O����)p�h0�����`(P0R��T=�"+1�.����m*~7z��Iɻ�0�":�
����!zT)X�[�fu�5�27��(�<ƶ@c���_o�=7���Yc_�A���B�o�|�C�XX��$5k����v�O���9�#���?��sc��g{>Rkĸw�$r9BMo3������0B,�}JBQ�L[U�%}��o$N�4\��"D����1%��B��҄�R7$ፒ��:�,�*\�-�	�ç,�x|�b�y3dcȲ>���qӭo�=���F��y�%E��x۝��K�kb����\�I�Aa�1=\�]��E�t0���Zӎݺ��	v$c}^��=5�`8��w�i���E�AKՔ:$�]�b��|W|v[�j��=����'_�JK