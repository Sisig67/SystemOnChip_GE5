��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��׶8۞�@�\ږwiܕÜ��=r(ro�fC�pr�L�O�q�;��?�����f��G��@�~w@��q����9-�:�D���lߙ��r�p�$w�
yf��׆*��`��]�*��Z����jI�m���0�p�/g�o��[$�(�� j~�[s�C�A/�5w�~�j�<ҷ�F���w+�ĳ#�itn�޲�g�rU(���MF i �0(.�f:�H�^)���|�l4�6�1�k�1�uk��)ckI+�W�����V�Y����dʨUY̏�!ix�C}���b��K��EY���qs���߸�:�.�I��c����_Ъ���d���d�pwfV��Gl��\�Џ�o<ݿ-dCʝ.rU�s�:D<�̋�u
,|�zc�>�}�F�5��7�{�Tm�E�՚p����@��GV��.U������V�
��J�Py�Տ��)KA͇Mt�ǼϏŦP�=�G�{r�J"Ɋ��W�Eՙ�t�d�9S������x;4.U�M$53$�_�X�5�q;���D��]���_ZB������`
������m�ä���)=��s��7�>��Y��o�+wm�2u��CF�1V�L�]u��%�Tc9S�=N� �l���A��v�b���1w�������L�G=��7b�"X*5)�q��P�%���4�6��gm}��0����=��\��k�w�̘O$�%93�c>$R�g����.6�׊���ָ��_��p{�fz)�*���>���?�y	P� 9|��1©�,��~b���&��$nVٞ�8NT|�L$g�e����.	�@m�*�	�nH��)9K��se�������>%N�����n���L�����B��Ed��?��c�&���vZզ8K���?R�&GF�4�'/���i�:qTA7k�0r��{��g�FҀ���ө~`5�2�\�]����j���2n�f����>Ak[�%�f<����%|�&z�de�	���K���p�̔�Z�����dM}���I;�&����Q�%|��V����0_,ֶ���U~pm��x_�Q�*�=򪝓m=އG��?�:����G��*�!	��ɲm��-.�� 6^�Lp<0�7���+ؽ����V����b����B����$�ފ~U�|�n�n�o5��0Խ�蛴i0���W&�h��E�k�f؛�A��v�V(����^�Nq��E��O��^Z=�9�-	�!�5b�3qc��s����v�S�zG���� I�����7C���pQ�V�	��C'��T��V���m$f�1��h�������z��/��aYB܈YB��.��0����y��凉,!2��R��H��+w�	�@~U�$$oK��Ɉr?e��.hO�����Y+����%`c������<sY}Tp�3���磎Y1�qIJ⟆.æ��Ǳy�n1b6Յ7��5q�U���8�B�'���	@'�O<Ԥ4�t,��X�ؚ���ؤ���G<�s���m�S�q��!��!@�O˝@\ѨO�5r�͈�8 �Mv���U��D��p���1�ЯbbBC�e��j�P<۠J�M��qN��*��K��=LffM�K��O�Ч7�#�.J=K+���J���Ҩ�M�$P1�=
�=�������tlo�ò��M6_�9Mrު��q�����[�};ܔ�*�*���h��7.[�Ӵ�lGoen�J�5 ȇz2�)Rd��j7!}�S���h���&7j�.�"!��,����7�X�F�ߨ77.���������Ę1����<$P=����=េ*|��a&���`N���&k/(���Xu���o1���D_��v��5�`C��&<������~���	v@����1i��V�A__P߼8!�X7��)	�����`2�A.��m��>zd9�>xh�6i~H|��0�HE�-3c]�����%e�k�a1��7+�\��j�iG�b��4*Oo][I�7ޣ��#z\YGk����6��{�]I�3�If���n�^K9��i�����JY 1�D,���ˇ�ԅ� ���!�:"4��Q�E��UT��in�	��`�3�j)(�d���/s�����0��2����2�=�s�⎴Ws���ԧ�3����h�譟��0@�7?����t��\�:�$/W�ho��-������xd��L�J,P��C~+���1;�:���j�-����t�2��8���jqHg����)Ք��?�͠