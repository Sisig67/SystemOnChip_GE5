��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���|���t�9?T�]'�=Ө��B.8��k�����F^yW#��������3�����W�\��U�mI5�#��A��K���A��]�A����?����:*�+!8j����rb�Mm�6��퟇�1��忥VD�,�*��sgI�%�1?���p�hP���8+DE+4��
*��i���� P[:_s��&O���b�������Fu8iZ��>��U3��G��'�2���nq��K�0��P�ou��UDneNNĒ`�'?2�6���Z��}jEt^jH�c�Po��E�NA?��X�̇9}Vf�]������1FRo�[�ch ��*��_�ҳ8� 0��퇛��Ò��PucLԽ����ԙ؂�{햋i��������5�2H$�,���JTѶ@�Zǲ�f���%��0�ޖ�'��F_�A��uf]Y Pq���3<wO���#x'������*�͎Eoa"�G����K�-�Ϲ��4����H�T:��	-N�Hn�M��GY���I�����T� ���A��+�e1�]E񹼷���M��Y��AU'v�b�l�kb�6�a�!G/AJR�xo1Ur;��N��p����&j�ibp�U�&)gP��[��9���zJY�-3}!��MT�Ev�δo(��e&���E�a���uC�E+�v�c1���g���"�YV�
�]|�.�c河Y��ݤ��Y���c23�����r��(��( ��-*���-������n�5]OC����3L0�G�]}�$�̥Uhb���oG.�:��vWAa�F:��S=�R��aە2<���	��N�^W�^H��t,����y�����2%ir�-)���#ʂ�$�k7;��ֿ�'���۬�v���_�ne���[Tm��jD	���?_l��7��T%���2��=ȝWrS��qY�u{�������?�7"�Ipo�H�����8,K��;�r]"��a����{Wk=H�-�R�+��nVJ�� ׅ�GE�@���TW�ѽgg�E�EދC(�����vx:/��r3��Χ�j��H5~_X� ��f��$��ܙ��gI7����4�:���w//�.�I�:��N����s�π:r�m���5�-䳣I��)Jי�>������H �T8лc�%RƢ��	��q�8������P1xpꕆoؗ6��ST��_s(�v������� ��L{� �sA=_���8�U�<$�*��&u/^!ܔ���yHy�6q�x�ʑ�����&"�5���Q�e���4��1_�+ �l��a��4R��x�+�7����4x2�ȕ�PT�_�M&�20���}bXr����Z�R��֛Bc��G �e<�XL(�?�}8��d�/V��l��Mg�l�R��P��q}/�*s8�D�;��fѼŗ�l�b,��XC�@�S�YӺ���GV\�/uW�
����+��Ԓg1͉�ǜ
�v��vt笖Phj�P�d�:�˦0�� ?: L���F�+j�'�3Y���A»� j��b{�@ԭFփ ���	���h�� �=&J`����,�����,�e��w����,}��P"�~,���R>�@��r+B�e�ZW�#�G}����2]�$%�\1�2������
v�Z$�Ї�	��EidI=9 ��Tr �u���g�Ӛ|�)j�������%�7���-�U��
�F1�	r*�"���1.����{i�mRUq6|�]��5�,�������?�"M�U:�J�rԟ4(�Qj��q�~�J��B$�o����A�5�j!>�T������;G;��߳�p��3�K��w�
�
&.�Q�+����>���\Hժl���ႅn�H�E�"�o��gq�[��j�:�ӱ_u�u�ЎSs���$G�����M-_4�))H8�H��Z�'��ZO���|��=ά|��u�W4W,?��٠K9��x�n�iiY�94ػml;~g�k">Wc�%J:��Y���e{F)�D�9�N�,��[�zG�9�P�-��\^!4����Ą� 'Ӣ+T$7٢g
��@����L?=�<Ź�G� ���D<�xU?9���	Fl�Q|N�rz?Pb�M㔨ǹ��F���>�������|��,���&�1u�4��Wc��ڬLV�cA/
��Ʉ�ϰ�ǀɡ�B��d!������iX�R�t�
I�ڟu+�Q�+�}��E��p?��c�G�,����y-�wvp���aݸ`��0̇͌��-L�m��n7 쮱�Q8��"��sŢ�-�9��	d�؏]%\_��(�#C:����N2�̟_����H&�&?�L�����.X�B���t���7���-\�RR�*���Xk@e%�=���d�Z��$	.���eJ��1���&x�7�����1�+��o��0���!qT��<ڤlMU,�][�pD��ɟ���3�Ԃ��A�v oH?�r��N��2BW������wn� �EF�؃m�OW���CP���u��7��`���+�������A�C�꺹>^�Wq}�`���o�7yGf`�b@Nz��.�x3��7��n���!v_��a�Y��
�����8�J��󬓝m:*��\��l��G�Mo%�thyVF�䘳�fb瞗0H�TigU��x��o��-���n���m�z�|u&`b��s6noMt�$�cJê�C��X3Cf)�H��e��ځJ�����$e���&)W���@#��fT��Tb�
	��]l+���^�1��R+qɋ�e������C�Y�K�Pa�ՊJyL�.d]KM�rH�I��(�}Zyp� ��1�>=���A-ټZwz�aӾ�xI��w?S���^�|������T��B���KՕ�g��3�9n��@�>�ο[��=�RN��ȝJܪV �,��5�*�d�9Lɪ��0������V��Q^L�L�SP�qݎ3�L�Ǖ���b�Ξw��x��w��$���\�>H���!��'h������Ӌ��{d��Ex֭^�^�sn��y&k� ��H|��ޕCݬ3Ň������[��^�'��+jv���Rc�?WFa$=-A�1���m�P��_ˡxM�䳟�`4�E� �����C�x�=�^�H��]hG`����"iG���E��y{��%�sG���HA�/�%��F ��)�fE߫�O�# �,�OGvp�}-8��W��j��F���7���9���x�����1��.����͙�Fpz尿�p��k{�w��q�[䲂'���C5�-p/�8ğ}���R+f뫊��PT��Y�k,[&S�y�T��t�Fy�&y�5y��-��e�)wu�NT�� ���_�31���&��n_�l�A���`f4���V�>B� �w�@>#�������d���	v�&�+<1C���^~�4��`y-��w��^({�za����h
��/��P
Ҧ�oq�%<��-��;FY��`l5$[���;���2�X�ڏ��W�(j�]e�q�ƍ��R�"��o�N�|ng#�����7ɭ~q7�y��ï�tp����D�xub���
,p��:�������Z���������#F�\*ξhfV~)kr6 ���E�[�X39��/&�$:��/=���X������}N�7bg*�|�mg�׈k}�Tg�HU�BT�ȧ��qV�Ox-(�{NV7�]�Hkt��\
� ��L2Y�6�+��7��>�7A��,X��.2��B���cG�53��3���dM�4!v�	Xe�c�tv|t �C�m� �T0�/��З�ޭ�̤�����*C_3*���|*Zd�fdi|���+6�/" ���N��G���4�I���pg� n�G�}Ă�ڐ&|��R`�0�M�����'�q�Y�pO�����!͇��gS̴���٠�b���������&15��3m'��:�ۡ�z���|2�r����H-���t��  =O��\�;�>��4� 5��X���wb3S�&'��ϵN��|!IQbAE.wFĽ��e�`�Z8o�Mh�UD�Z@Ie��;�՝������.���ң���Y���T~8���Lܹ�-��7e��m����g�d���I���w�[��P��#D㩏S*������<�<�cQ4Gk,&2>�����6>��*��O�"�Bk;)SE������\��q%�uh9^��Կ14�#lM��D�˦��	��)�l������T�^�&��h�Z>@���%��u�_��ʜ�/�O�yE�m���X�t
��L;�N���\��[��0}�oz�2
݂ԃ0?���G���B&�;�	!�<�G�ۓm�(���3Â�T�xe ^R
*S���R�4���,�aO�7��_���tk�J��x����.�D��m���G7��T�������9�~�N�a{6(�_����G
� �d{�f�0��sh��-Y��O���f���iV	�-]�H��#a�7�dJmo���yL�c�땼C�l�g���ͅtQ�0؎�a!堒�'K�d��� ���(ۊ�c ��(Վ�V?�BR�'�cYd��Y�J�:C5�tJ�2�=��@vRP�0e�����ݑ���<Ks{<p�#�?���,8���-��'�l���rQ�)_X1Q.��j8k��p�%`��Qs^_�W�L�E��ъ��]m���Iy'c �_,� �&���t2���lST�D���u�*��lj'1�짩��3Z*-|�f��_�����1�@n̰��̅�#G�kae�����w�%~�kC�i>2��<:?�k��Ib��(�Q՜�㼫��Z'WJ���r�m��K��w��-�%D;^|A�LX_FZ"�9~;��xg��g|�a���/P����
�:�����,���Ͼ!�7��)^jǩC���}5r��ҴR],�D�U[^���f �f��ͽ#���� <�"p젲��т����-h�c'i��=��_~�7�Cz���_F�\TuF��m;�F��-�
Y��7"���${c@^��W�r�/�QL X�� ��|�,�=Q�2gA4$%^����i`h+�'#߹�5Z��k�é��H�d�c���D�_����?R�1 dX3?�˩}�r�MC'p�����"��#�k<���@�0�ٮM�8U$F�%Fu�c+gA�	�M��4=�F�x�8n�r�`(���e.S�$!�A8A]��xy��E�$g�h�V��Չu�a�Ǡ�� Sq�
r&�LV���w�N֠��o}j�? ٺhz}�Λ�����!"��{H�ٵ	�Td�'B��mӸ��]�w�a�8L�-?
�'b*����dQr�g*M`�Bә�F�����Y���ɏ3p,��Qx�ݷ0���V�TGC��(ݢu��ǋ��$�[Z9��{�=UX�:���%�4�{cY�^���Ԣ=d"yH�����S��ڃ��cSi���0F!���P�Ɯ���`:��8ܲt��ѷ�}�b=_ �G�;Wϵ��O���n�	8o���r�k�gM���E"[�EF�[YI���3�a�)s?ܔ�t��w�H�Ӂ�fwb�N>PTL�NMOW�I��
E9�w
����("�PмK��|�%<"�D����ٍbB�j��X�Y�����Gw?!9�'�ǒ��;�D`�x�]_W��
VӶڶ�G0�����Z�L�ەd	��N�{�fL�'��n�O��\2�rW�eJZ;�z�/S�va¤�Wt���=���U�Z���7��H/���Lأ%�@ WZ�f_i �E?��E�ьL'���1��`��υD��5A�H�9LN���^�����8�3�7���S�ۨ�G�#F2�e�Uv��-1�v��X��vl?2ce�y�NA���9����������E��뉷��݌Q
�#���wj������ֳZ.����Tm��	6�^���Fk��,�͒�x�c����T^���YSB;m��>�A =�c�o��o����^J�*,-��/ԩ4Kiz>��R�;i��Y6Rz�J#`kj����S3�Z*�\xI�)�>f���:Z�
�������싢0�oעk��	���m[u��f��،�y���qE#$i����H
= d��VvM�wɖw��m��h�&J�� S	Y?�Pی#>�
���*��F/�����!/CEz����%� xx��%S�0��nSS�l�ﵿ�3�wzT�l�	7�x�[B�~����Hǟ��ji�d��ώY���}��.�zX��X,j~���(�����a�yim�C#���}���h�v���Ӛڥƿ�d�5���h$������c��)_��y#V��3��"r�Cj�K+�^I�Fer3��I�?t�㫽^�2�sDP����Ї�:�1H���w"�}�� 5�G�_)�ihhϥ��R��&7"�}g2��xP���Y�WI������Z�:�p>	&�f�`��X���e�E?�a�Wm#ױ�$oC^��ޅ�����l���"�٦S龠�(a	׬qdv����E��O��������T���1��l���D&<r���<M��H��3�Rg�)͓�k�y�=)��T�>��؄-���t@/ӧ]�4�E,�z�K�a�%'�Tn��S��k��w�:�=��M)ڻ���x)}P�x���U3�ʅ5�|�����\���. �#��	����T��p��s]ݿZ�R92��P��/��!2���<�O+ۋ�t�q0�Np�w9AJҚO�LT@����i�~�-2�(�J痳���>U��,>Zd�5@D�v!\��/��Ǔ���@�����k<�'(CU;\{��f��9'��I؅�|�[P�?bp�0��Tnt�
5Y�����	��y�)�^Ê@j�AV���8�4V)�¢���s%S�7��4���fq�G`�@�tō��ҳ��J_uV���`��n�H�{�"SL��+�|��ㇵ!C��L]/��;�/"��A�>6��yޓRn���f��7s.���H��kP��r�cM����3^u�F�{��NGN��3̯�-m�B��L?K^1p��I� PI�>ou��;�_�J��ɬ.� #�0LrF�ڵ���_q�r�w�� W\L-�ۣkC�%��*�����ː[���%?K�M}����[w���7 �a��z�W~��z~� �B�9����E�|�$�5DM��b`����C�� 7��~8J��T��xm�����Ѧ\��6�=���\G�3p�����������ly)>�iӶ?E��Q���J�`�/˞�D1��7�PŮ��:��n��l_���z$�X����I��;�hz`���e���n$5!U��Jq0�~5ٚƇ��m�J?ۜ��)9D�&���'N&���S�X�3�+*�2���>
.�$���H�҆/��.I�V-�.���sʖ��� �ǓF���������yQ��x��;S;�c�*r4?���`ĩ�)P��.(!-�압���K2��V؉���;Ε��E��C� �V�&��S�%oQ���%g%3�N"�6@���~y�M&qU��,/�`2=
�ҿ)9���`$���p�����9m����ea�;Fd��=�&�+�JyY�xt��� 1�`���*^�|y��� �.�h$��O֤�L�X�3��|��6���	�}Z}T]������$�?� $U6G?L���8�d�6�DA�Yp�۬�V������{�$�c�G����OZC�1̒Q,I�b�qv_;u��x&�غ~��=bА`�r[Ͳc�̎�W����}p�W�K.~�g��7�V⸇&�V�s� M��1׽8b��|�����Ѕ���+�ϯ?�,Y]t͍�����\�_��F*�|((���c�#��u�Ipϲ���HlDᑣ��	'���(���3_�Zc�Om8ՙ�'���\f)x��M�f��u@�Yy%�O�|��,��sh0����n�Aذ/9��K���ܔ�� *m��a"���0#�s&.���S�G�M�:�t�N�z�/�+������>�+#�׼m�i-]E���N<�d	��T��c��l�_`}���:.���Z�z�K�j�l:(R��z!�'��>@��@`��Y��ErgCC�r�<�-���6��տ@=���?ZY��bС2�ߋl?�:!]H����.�Qu���Yt��ȋ#lS��_eB� �U��mA
2l��_�G�(m|��
m�QϗM�@FV���� aH�O-�\7/5 �Ge��6[��w��b��ᢽL���,1�4D{%�욵��[�A�&��~��A&�=r������,*4�ͲIW��c�f��oy�?��n�8m�2�Q=�.�gba
ˢh$%��ޅ26Fвz�4��w�b��Y�D\�wI��Q�T}�O�>}��םc����a��h���m<�½1j�������a]|D^����n/���7yMI��V�o�c��w�Q�������5�C��<�ޯ�pY���I�G�\��鄅�ĵ�/�m1b�ey����;���GPS0�N��`�q�|�>n1�JI�����5�h�^:�I��o���c�xӔ�����oP���c����f����s�E[V30��{.7c,����e�i�2��H}�R`�v��A;�aя���Oz���b�4��e�E�폋U���S�5b�\ZL�s����[m�T��a��&t𸚛݉�r�2�%#Ye�����l��n�U!��c!��.bv��5*���n�	I��Hp�m�PDk������+u���-�[+I�LpOb�b���EO�(�O�o?)�go�)��-�c|�EKwlkO�PVd$v�{ik<[�nȼ�1�1�p�hĚH�;���׆F����ͿH~��1[Z���`z�BP�e�r&�ʱN�\kC���ء�9�2�@F�[�踵+�Ɔ�f���Y�\<�oN�\��|�3z�5<��?N��K%Y��&�#����FxN�H��0P`��]�|��8؈�i� �@39���z���\�;�"|ѸbY��O1;:���O����#&��;a7����4b���Z�i������R�00y�<XU ��$,=&U\\&zK��p4$zS�Z��� ���[)y��r��:I���%���Ah�8�:uP9�������g��Z~��m(i�	m��E�������qc��p	�1�1ʓF�m�5sjoS�V��=�w?j�2y��<��o$��Z�+�V'�U�u�%p+X��i���>˙Xjt]���l6هF�ٶ��u�yGM�5GBw&-#|�b�K<�V��5���j�ܙ��y�������PF�MO0X}A�e�<f=�R���ٲ>��@1��U�$.q+ilm�q�]��:��ќU?�<r5/S��Hȿ:��H\WQ�,�:��2�H��3�y�fWtQ獢Lm�\�^C*�@�HWt