��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj�N���0��tK� �Ī2�r��$��D��P9�Ơ� 8�H�9_�Z\�'���=n�?�r��'��<�I��"�Ȃ8�v��s�h{<�lx��̄���ֵ���"}!A��k/$%��h�����
�aݲ����~BԄ����$��^Cr<�iC������T�k.�\0/�!���Z��V��0!ܡ/�-�ŉ�^u]h��b�'(��ϟ%��Ł�Α*:�:��L�Ր�K�a��qPm��R�����N���J��zt4��B14�����7�܁B��^��\�ƴ�;M��,N~b���X3q�n����pb�x�Y� ��$���
�'
���uaܗ�WIg4_�Zd	B+�fʋ k�[#A���2f&p/���󦗲��jA�� 7x��lh&�ȥv{_+��'
sD 0ċ�*i���T�q*̱����:�����č���3IG�Om�ô��Pu�J?"�@��K���T�N��f�2�Gv���+����&����;=�TTߺAd)%��t&�R	���RC.��H0��:lT��MP��}��~?����@4>>l�ow�C���@.��r�k2�@���&�_�ܵ+��)�oђ�PP��8?V򍂵�9
W��l�ש:�vR,��tNpנ�1��ײ�5ΪO�*�l9%�9�Z��4�v��'�5��Do�w9��{���j����߼�R���Ӝ���ٙ��E8�5$ީZ�X��Oŝ�#Md��K�G����@��|P��U�=�F�2�����ȷLe_����.�R���QF��A��!�Rr�	�3����D����$.���!��WT�A��8b�����h�����$��(����Ʃ|Ӹ����ڶ���]i��Z���>�w|��ڀKk_x�O���������f(Ph#��^��iI�J
T���9bQ�2%�簴��x��t����W|�|��~n��Q�<���rҁ�f�����^:p�]Wu�=���� �F�Kw����$n��}52�VNf��}\71�X�g���:��"�n���3�ͪ��p���Y3M��H���;M�r���[�a�`3XM����+<�S�OrݬH�6�� �%�g���
-�mSVx#���~�<"_���HIz>��#Z��&�F_o�iI��O��)]���=�W��g������L�.c���J�.��}<4�?^K\�Ş$mD�r��h�I#~��= ��5��3K��žl�.�T>���tË�kI�7뢑m�_Kq�c�y�mlr$]����jپ�K���t@'�kO���� &��IU�L:��t�K�5�����r?�~4��e�Y��w�o���=ܾ�29�Օe"w�V�xo�&��s��]4�<����S`Fd�>.װD��gɛ+"�M�js	�pg!ޢS-���C>�Dng{~T\�E��*�����i���;}�M�2��M3�
�cWS�H����;A-1�9p�@��AK��"9XHs�^�* a�#�is�`%p�C�	��_�t+������2�Qx�e�L����j� ��!��N�G�u��i��}o��p%��؝�E���Mm�[�����D��A>�G^)��ǜ�^�x�������<��;�:�u%��Yu��C� 35�ĳ��s�;��?$g'��֡�>�5�X9PLF�3�� %��|=�A�$xwX8'��~������W��
H��P\�ٓ���|�Ry�gt����}��A�|c� Y%��"����n3Ɉ>+�C��ݰ��L��I�dB����!��[��ڢ��$ y�/����e�D�n���0{!�!�;�lf�T��E�29�/�{�D���([��U.��'�Sl*���|#�?	���z}V�H�ծ�Dڷτ�H�*)��B#󁳷�C�^��N�Q��C��8�}%vh0���~�A�V�k�(g�q<��/,���Qb�޲���곑���ۆE�(�H}T�i�P��q�U/�"6�{�JB��t)g,M��!1u��YX�b���o1����W*��J?�B�Oc�"TARMǕyϨ�.Pz?�
���쥻%`�V���Ǆl���,2�*}�2c����7���j�TU��X~���oH�u�����?l8�q��������c[Y�j��ᇤZ�=���5�O.,�!�
��70kF(2BoJ:�^���+�ßA����pV44���ؗ3w�S�:�:2I�ܬy��h��!��u�'�������7�&8���R�^y������J�>�jH�GX{�S>�J	�ԢAf_�ܕR�C�|�%���,O&�t&L�����J)�F�+���fzw�6	7��a5���H���
��u, QK��R�V_�c��nM����]&tLl�����qwZ����!qim����I�S=�{��,��1I�z�_F)0���$��AG�Ϲ f���\+b_5�-Up�����+w���s�D��R�
�k����5�m�:/�`:�/3f�_2�%X>t^R�����:7Z�Wd?��J��f� ����u��_�x��g]#]q�V��*�"Ǉ2!��Z�NK����O�^-��)U�ؘT-"L^��F��z�L�d����\��6u7	�2[�T��!X�>�J���
#	��2{`ʓ��"`��D��st����x�|�_���a����AݮEѶ:��{�C����n�O}����Y�]�\�O�X�[�e�KX1���R.�v����H�V����ݒ����
�&eȱ���a����w+S
�����!K£C�FQ6Ef8����S9Z���&�h�gK��:�0��$���B�U�F $D�5! �BgϷ-Px7��</u[�*��;�I����/���[�i��C���#.���L ªјMr08y�3O.�2MZ�J��R����E��,o����.�b�G5pU?fLo
FۚQ��>9ۦ��N�	ٯט�z��Ѻ����H��lZ�S��$UF<}�eQ�<ˋy*4���������<2e-
Z����IEq����ԃ@��F�gb��� �@�����Z�P�ēNYܳa����a���s�I]�?~������e������-�z�w�3��:��OK��O8�pB��^�吚�/G���@ ;����٠u���-l�v�'�-?C��J�����������E�~��Ls\8i=I��9b7��&`8��㒡�uP��ι�NPn�'��$��p����o�sJ�h�:� ۯ=����%��呇�r��Ŝ�@n�9A/c�^�P��Y���DNT��S�8&_[O+��ڬ�XKs#_,$34�?���{�|�k������\oQ��VF�o��T+���BcP�S���jUh�G��ea<��ͽ)��<�`�3'S�m�ͽM'�A�.!zz�A�}� y�*o�����c� �@jd%�4.=�BK7/j��z���XD;�J'fM�= s��X=��)�<<'2?�ݫ���b�^S��D�&��;	|sc:�%E��R �]/	��9�A&��#y�q�@c�ø���Iw��)�XS�4{�w�k�<�+��#Rg��8%t\l���W]�l�s���>N��ZN�B�C/#|��.�x��WR�^�E}w�Eb�W�K�'� ��(;��-�M��\lb.>腪@��a���t�q�,�l�ym����?��u���:��V��}�!����]�傐Ā�0����������8�+zd*�ބ�\�=�N뭢����*6�����<]��0g���|�k�b%��(_����$)����S�t� ������,�ݙ�9ާ|��<ˬ�pS٫	eSӞo���y>�W$�ώ�5 ;�F���)K�Ѯy>s�ܧ頀�Z���`�c��ܷc9H.�������$�������T6%r���5A�lu������m�֏�'F�ߒ9���t�Yu��~���A�X2b�V�@���
5/���Pq�$��{�0�j���9�K��Б���}��