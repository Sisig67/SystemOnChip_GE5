��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%��%PU�>�Ӱ�~R��<O��H�I=D������;<��y~O�d��$�y��y	��L|��]v������p
�)�M��X�_i����d��mm%���.�Ð�7-�MslW��p��AMm���k��6]�N��	J��<㖃Q�u�/-��h��_��D�7b������2������"���T�>p]��T2~��B	���cʉ йY�EqYf�4b\��+u��q�!���0 ��¼���2�_vʟWn�X�O���Xk��m��h����4-g`^���9n����;lݽL<��A�%�����#n��]����|ޯ��gYet^�z)�$��9�ǝ�\6��]s��J]�I7�8��||�G�<P	��8���/v(�c.��l�K�4�Q�V�턿u&^���b���m�����2V<��V�i���j���"���A��gf�"*Eh��_�CGU��a����	�l���,�#u^j�dcM�Ӷ32�D�)�uRY��F��A ��j��v�9Ѣ���'!��f��/����-������g���oɍ#���n�9�/�3+:W�4�M��_���p���h/>=	�X=D�sq.��gR��ڵ'�(��z�B��cK�v�A����ߚ`l����3��I��:F��D����ح�LENm��|�B��?�dD�$�\�8i���~)�`��[�I����(�]��R��L�0X�Y,uv�s�.膯��#"9���~�:QTi ��߁5�a"�H�.���PP�ӌ��hK��f�"��/���^�J��PG�^��t�YV�3�n�ЉY���d���^�k�z2�,}�q�2ѨuU���V���<7'�H'}/E��i������H���< ~շ��䣰֐����k3@��� 3���=d������/,�����.e@:S����GK(}�ti���\�j�^�b
8b��
U����`�@j*oa�ә���j��˨I&b<;}Gn
׻�fm`\���Ҵߐ���`o�B�HZV���l�7�D�3/���ʘ�I\�#=+������8���4���{9��]p4���.�C��O;�$.l�t��@ E�D��"D0�T�7C�n4$P<5*��{��"tKq��M	�� �� ���{�;��z'�G�n�T�˷�
�=
���+�3��N��	�{vI����*0N��S�gк���0A�A��}�SI�t�q�3-�f-o|>0Zld҈�5P�o�����+���&2/���=�Gh��rvy�����Ex"�%�~\m��q����(�r�q�pX�� �L3\O��3�� ���:P?�.�2���py��H���j�(Q+�%O�\7A9�TQ6�a��f�#Vr���9U���}��Pr�*Ƽ.�|<ݭ��"O'�t(f����r��v�&j�����	�8_�[���~�7����!�5�qcF{�k�`\S�Оﹺ�WBw��� ��3�zJVg��|n����rK6Cj^v��1�;�Ok��Pps��h�K�!�{�s�Jb�@Ii]m?h�4[����Z����/�)Q/Xߊ�*������nR�}z�bJ�Xo������/�Z�^JP��{r�O�`�f�r�5<"E����k��Z&�'��N L�e}�tf"��5���[ő�3�tiף�4(���8s=��al8�$�;��8�;�%�N��)�����:^�� U��~��N��(`ȩ��Ԃ�z�nI��hB'<w��Dɼ9FY�M�,��H�>��7��ũ���8�|��������n�_����\rD���I=����o��8��D�\OOB���I9�{��h/�@�0n�IƢ�fܐ�n�X�\�N��F���_�7��
��KwX9&��>~���[��L�iW1('��/�Gt�~]Ys�5,O����G��=F	%�:���[dO�R����zE�`��|�ʳ:�'�p����`o=��������O���7���V�� ����cL�_:��8ݵs�w��^2�x�� �Äj䨑�t?��� �ڶ�-O��̮�<Z�}<U�����ƙ(�۪��DѴN�D��2?J��3"7Yq�}�|*�
=*��H?@�F��c�2M��6��͋Q��6&g��CEy�?�7��-��kU!ť��~e
�JL�����A"ݢ|�1w[�CÙ��u~5�s=X�������q��|8w���]�D�{]� {MNM�+�"E�7�n��|��G�����y�.�?8��*?ov�$�d�vLj,��Mn�	L:y�C=��=��g�g��������(�+dwB�sB��&u�f�ձ�$+s����_a����5?����ihՇ-*�,�#����,Rv:��a:һ��<�d� ~l��K�������r)M���Z(�����_�+��C3�:i�2z���LY��I?Ao܅�b^���	h�p���s�T�x�n�r	�1�}!s]��U����x/��3됄$���mMi�+��)��0J�ֆ��~�e��A�D����hTV�l��(�yV��E�jN�f�뻍S�.R���o����61��������MzQ,�Z���C��f:�R��u�yc��(�&�*�f�w�Q��a���P��w�+��f��M�N��^��1���rȓDbDk���0.��/��)�~Wx^�b�AOQ�Lfk����|1�oy�D�������q�ܠNG*�u&�͖&^��[Q��u�ѽ.(���	/���&���G��k��I�˹۞�,K���ѣ�D���;�#m�c#�H�v�(���+�$�9�֋Y�����H�f��C=�;�`W�tO���칃5�G)��7�ǹ�����5
��t����Io����!t���A�W	����-��!����$A�Y4K�
$���%Q8�7������~��I�_��{���w���V�Z�(W$	�Z�"w,��B���h��bI��y9�
��a ��Y����x�E*ouT��Tl#v��#z�~�)Z�M��\�����|���h�	6����?L?X ����BضPCd��^YX��7��� ����3V�o�t���R}��ׄ�6�.�Kr�sN�E��hV�6�X1i�,�CF�{n��\�z�Y���z &�5s�uzWnv��{�� ���n� ڡcN� ���/j���,�8�z�Θ�A��x���Ƈ}��\Kѡ�+����������b|4���]'������ط��S��-�yK�+ɓ�����=G2�*�̋����p�&V[�~x������/):�bP[�b��P8٤>,��C=�B����fO�T|�} Dk�#_;�>8��I{`�+8�t��b�Gb4N-3jO�jz�.����\��bW!�*�yc;0������k(K=m����iHo����p�HؑЁ8�Gs~Y���^�6���\�Tlts��&��Z����5��4f�1����ǧ+~��|� ����Uyѳ�\P����Y��]��3��?�	�3d�{-�����]7<?cQ���'P��4��ݝO�Ff]�;i�Ņ�0�]�.�/�;p/�̅&S�Y�`�Y�3�f�����j�����^�cJ�s
:.����S��a(�ڱ�#6��=^y������ZJ�>��w"&�@H�=��`N�Vޱ{��	�ؘ�X�ѭH����G.Wih*qs���ϓ���2wp��v�~~�i�
�9���_�s�f��d��:ݥ|�Q��UF�����,wr�
q�n�hg���F�	��H� �p 3���
 �*��%<������v/�^��ps�z%�2{���{<��l��hG����Tr�!P� � 9$gmY����z*�v��P�H~VnN�_,�����ED�¤��1:�s^0��i5	;82��z�PM��$��!�^���p�
�(R��ȸ�l�C~�=l���#W5�tϲ��c�C�w��5=�{��+Z��������9��1�����>(ǜ���M)����9��Cv��-cd��Dk����n�{Z�YZ|�b�w@:Q�\z�>�0����V������|��q�T��-m���%Gk��Uc����z�Jـ�D�p�Cv�$�������/òq�;c��qfr�:?|[��@������*�I=��	(����p�������T��5*Q�=���Pï0����&0��	Hee��[��o<AW���#����w��[E�n���8(̨��>K1J��}����<���;uu6�=B=���zo[E���'WBCM���'��K�Z4n�"&w#Z�4q�W4��{B�E���S��/9I�`4zS����v�Km��%sJ�����A?pD�_�K�`�/��#tk
�q�S��s���6� �#�5 ���Z>���=�5�"�Π.>�d�'����<+|	{���޷-#�O�����.��^Ժ���_脷w��RŎ:�ԶnAC�Wk�/���+Ac��m��\�`�#�a�H={�$x+�'���p�{^Y�
�د�h<��ڋ��]�v��(�����Ÿu�f�̈����X�#ZU ��8!�}q��Q4o�a �[�h�?޶��n�{�����2��䣊X�G}+��>�T^��3*��"�h~�G��tP�� J�&���F'����n�
q����jV&U��ڈ囦�����4h�F$��Ӿ3�:ln���['�~zy�E�_�Кa�����sqӾ�l ���"��:��$r�4<&��4W�H�8�YO�F`4�.��H�z"�u�+ߩ��5�mLH%�W��D\�c:8�UW����Zs�~N7Pg�B޾
%>���n��|��IQ�ގ�^��g�О�����P4_���\��H?`���0�y�~��PI�UD�m�j.5�7c��Wؑ��*\�Ma=}�(�)�2��}�>�X���S�䝨�m��R�x�[V�.�N�0�B��4f�ü+�����h�((1 ��5Ձ��_�/�X4(�p֭X�u��,�ˈu5�僾=�y�g ���K���# őB�I�/�Rm.5�dt�<b*T�(�����f���3��G�J�	enc� ����7� �m�^tt�|puM*�6S=��iZ�%K��&!!	�׃`ǲ&-h]����<ݸ�D����b-9�.5��nIQ�t���M��u�춼a�>V������Rbmj��T��;�JĞG�eW4�]�l$�利5�U��S�`��y���'�J���a��?4/Ԅ~$D�4=�$�zzT<k1+�?nR �A�v���θ�☨x�WSa�9��r$�!yS��F��%c@��o�n�'#�s�qG�DRkN�����9��x�ֲ��SA�D��n���q��o�����tW�i�F~�!�5�^�cجnĢ	#����ۃ{A*�U��]ޥ~sܘ�$��%Ws��FI�>�z���wUm�&�Z���1.L� ���=�}� j����4ȃ�\G�|�
YY�� �E@	��Q{�.�r^��2K��zwӨ�A�~g���Beڔ�U�!�#b���B�q$=�.x����>TV�72���v���d}�7b6���ÓT�>��TO-s���-��ߗ���X�)u�8�C����FSSj�}�(��̖�?�� �X��g_ akYʉ{xq���}{Bx����B=�o�^q*ͱ����U���ouR?e��F��{;�g��#;�3冀�tF�jM�ީ�_��Ȧ��$6K��ㆊ��a��Sǔ-E�x2����l�I�UF�}��4uѫ��%��\�2r�O�%��,u�x+�b������&O��t>�N�,cR��PE����N���GN���*	y��0皿��;1��i��ݥZ(��4/�$u�����ȴ "��B��Y�ؒF������$�Y�4jC�����-vכ���e�������ʢzl�'k~�݇�u	 S��֐v��h����m�a��<�7&�;;�r�) p? �B�<"Bn[�bMO�Iʂ4�$7��O��&z|�����s��(B�(�� �*g�&PIj�8�2��8��I��0�1��'y/eݟs$_��N�z�?Yn�3�r��{�&X�%�� (�\���m5+M���"s��BBWk�� �I���[%s�v_���˄�,n�v�0\@6f�J`
�PRk��&��Rs�I�k=zR�v���D�mFG'��jb���)�*п��fȎؒ�HI6��dr��߈�󞥤Q��/Z�Ν�#n,iX]e�>_�tUp�?zo�e��U���Ak�؁�ܷ�gV�l�����v���鏆cI�KOА�\/�T�670%�Nr�ȿ��DiX�x��ט��!�0_mF�0���X����:�=�7���i8�?���ٴo9�5�����rӃ�Ǐȓ���U(xJ��>�6�>���.���E#VEe�QR�����m%8�N78��i.kL*�V�?Ӽ�O�G�o�e�U�¼O��WB�e71�|�F4%'u�ɕ��	���5P�@d�H��o��{�7Hwh%� DŰ�Du��R�J�$C�~�����X��`�0R��_�����\��Ϡ�@�v� �ȁw��+��@�[=�bf@ǧ�T��s�������gx@8֖�T���6�H�-�����ǄO�<���8|����ŁM�3̷g�u`����Za�Fr����47�XX!�c��2x>y�{�Bw!9�����F(����t�M�#�������WUR1�{�$RG��9*n���/��η�5fc),~F�4o����y� �團K�-_D��{��frS�H�)���&R��0q���z0�⥽O�e.��0o:����m����1��ߊH=m#�u�cH�P���?��.�j���ϰ���n ��7�te��yA7ڴ*ײ�ܠ*��0��ce2X5��Β�d��$�!?�q��C�Y莎|]��_�	:�`N��ٹ��Grx�I�}G�+�������:d��{^������8bMQ0���l��>'�����`�r� �P*����2b�ek���.i�_��������R^��Y4�I�=�Ϋԫ�迭�p�5@X�����\�g�e�g�9���T.շL̏�����#&�j>*3c9!@tL\j4װzT}q��3؀z5ybld(a'��V18���8r�$!������ӽ'ʭ��������48\џ#��5����/����afGh=����nx��6���)��;�>[NzH;�P�>�;H�ʺDM~���(�5Ȥ��1�Sm� O��Er��iP�@D����9�!���\?��
F�/y�PӾauc�8%4C��Q�u��������qB+��Ȗ�烈+Kg)`VZ^g�  o)�έڮb���[�8|f徻a¥���@�lCER�����������/�k7o��H����HaQgvS<+�}b����u������^�(�xUq}�"�hu�jEQbJ:�a9���)��9;����:FHY�]�t�¦U������Ur��*�Kɮ?�?�w�6|���VTc�Ad/���Z�d9c�Ud`(�i5�p
�\T'�`�FH��'/x����e����(��ƁĴ|��j�h���,.Q�hޅEwJd)�	��^d	��Sn�$V(�"5��x,J/2�X�1�ύUWM��}2hr��Ǧ���z%�^Q�$+��Տ.�J_cu��7�����Iy��ƣʗπ�1O&{[ �e���D��r��qsv��_�Y������� ����K�S�cEo�~�5���X+��K����)�F�:�7�p˒cta�������;���*��Cu����.�p��O�i�{��ԍ_1̜R�-�R��=.��=F�"G[�fl9�����Sꆜ<�6�ǌ{������OJ���c��yX'�'�[Sߌ��비ۡS(���g\~�����l�� ,��7t�	�K1{�n��XZ֑҈!���C6
:��.7�.�W�K��=~��Y$�N����(t�W"�ҿ��[��������J�ƽ�@A��؛���)̄7u���^e���Q�xl7-�����FDV���J�
"�7Z���J�)O��:<��vP����Ȧ*�md���I�SӝѦ|��r������Q��Ρ���-�~!��1J�&rp�,���Ν�y�'V��jpA�*��7���74��jֺMI�R���x��ï'���+����)f�R�a+�J�g�V��O��s(�aH��Z�E���|�H^!Fj4���Z=�i�0r�5�h��äúti�y*&ڋ�!a��.�i�*�]��f�f��ʉ�2i�Z&>�v ��|���Ʌq���A��w�g��!�����-���G��܅�Bn�%{�Ty΄�c����iN��.F!N�I�"%AS�M#��� ����T깵ZY$\�[�$;m��qs�r�d�K���H��F��G�{�y%������v�!�Q�A:B��h���K���E��U�2�mT������G|�Od��
RU�H����5�7{��4�Y��4%�PH�*��h�8j=܏���Y-�qZ�8���rIO$�1U�a��n�A�Հ�ƁSd�,Z�f>1��/��#",�ؙ�V�~�T>�Mٶ��XQ=b�O^�Z]9��՘7Y�d�n�-�WQg��cD�=H�Qk^�I�/�m�����ϢB�#h/N�bJ�B��8�86��n#�o�C冂a�c$�@��U�$�9E ���!Q�,H싍�B$��z�Eu�����&��d��H����I�'���6٢���t$�qc��� r-�r7G��Y3c�q2�a���5%�H�L���IOm��h��P�g�ϣZh)���ɚ;B�x��-ּ���-�[n�d3��}AU@��F��'t��]Lf�z���Jʃ���v��h��+���:k0]�*^T�i��0���8Kpl�@�u�m7���P@�'�<�$��	���A��;e{ܣ�m�$�S��o8}@�N,`���TpOM_F��W�N�B���"��ǹ��A$)d���A�Ʀl#zS\�|v��O���2%��S��B��Lg�&���æ��a�N��L����٤�S\h4u�w����n�7R�s����K���3"HZ�*V(�I��ڷ�(=%�I&tɴ�kR����a���ۼثi�����}[Xڦ.���&s��T��tѤc����2�Uݚ����K���BYy?�.���d�01�~�B�5���e�[�ՔzxK>soJ_���eK� zS�sA�:ZҍSPe&�b_�q5��
�,� %{h1(<8Nʴ��t �Gj���lM�u�9��5/8(��6M~�:�5�K�+�ǚ�ּ҅��U���E��+��2P�>�1|�Q�|yQ�@4o,,��z_>�O<���&�4�l{.ibj�p��Aά�z�f��!>R;�;޿�D�E�RW')=�dyh�HL�I��{.���3�Ox�N4N~q��Y3���$!���X �AI�Ir�͢Fp9�!�ʔ>/LC�k�F��	S, �T,3��h$�b������X���m��o�1=�}��c��H���\�-5���C�.�����4f�횵ۦV�lRn���ymr�+��ե�`7r^i�j�
�1��.i=<��Y ��bǣ鍫���dbt�bC�2��˶ޘ�G^:��ի!�����Y:����M;�� ���?h��7�SE5+7����4c�.�B���p�x��nȽq��QA�t' (�,e�?�4E%yG�u�*h��)#T���X��^���)��j���M��=@X�H���و����E�g<¬9���D������C��F(w�qAܨ�3c��@�j.��c=���K��ob;�LV�_Z�gtX���vq�K"�l5�7��
��� ���}���\�\9rs�O{c��'D����ȕ��`�5rF|�K��v02E��%�t�}�5C��E�
�%�Z���1�^���'�'ʦ	rO@)��)J("Q�I��2�n�9*ѯk-��x孥� ��,/ҽw[���aSMl����an�~�%� ��h~4�
ON~�n_ߒjz�ߒ갂ڢ���PPd3T�ʼ�LL��Bt?5#Er���,Px���8|��+�n�k�^&��#����˱�j)�H�J\����: wHKr��C��a��{�ě�0FH@��g%`���x�tc)a�z]�6"M��ѣj�l����>�Ff0��y]In��`�o�G,�#����?��]0����`Ϯ�_~�y�!�\�>�Ծg ��I�D�0��K��l��=6yݦl��]9��)������1XN^`��a��񹦦Se4Ԟ�������$d@�n�taX�FR���ȹi�`�C<���2��{#�/'F�E�H$Sm1�Pf&nl�-T��G9����ٛ�]h�(^�F�/� ¯Cԑg���+���T�2�		*��z��I/ɯI�h�?�N%y�G��Z�O�%U�6����
E:�mF0�x��8�oN���:�S�޹"�6B0%#��/hx%e�F�i�X{��*���Ľ|S5o��<xS?M�E 8�|n��O�/VpK����RVk#e���֊;�����&q��Y9����F܇�,M}� ��7��`%�qi��f��&�sp&��:9\��8���{�>�_�n_�lKocC��8��s4|�4oݓ�j��-a�4}騻0[�h!��z��\���r���8��[�wNuF�^�~�2�ˉ9�U7
�
��*��f%9�|S��vۻ����8x?0ŕ��G�ϱ��2)̔���$��۝�~��")mE�K����=+�1�2����qo
�i_Q����� �6Y��@��I�]"�(���&�C�'�ǆ�Y�_[Sq�_���hGVn�̱�G�� -
�-ӆ�b1[3��:�W�p��G�(��ł�Gȸ�#�:4��K�פ-h�ޜ`�{-�-7�ʚ�x��%&���P��6\K�a�s�>�PC3n�/��Y�]�TU�jdhv��W����K�;E���V�0�a5k<�ѐP)�,��N�u���^q�$����}��<9-�{�3PƲ���k�7NH�L>:f�3�	�డ9Ew��+�|A�WA���oݑ���e����Lw	j"����KH>ƥ����@T\,���{F��8�/ņ�£��7���Di���.�1�h'�Y���S;s��:�5�|�Q1e�~cNh�Dp쩿qOp��m��L���6�IͿ9-���П%��B�oP�׷g
Kg����hsf����I0�g��|0I;����t�y1�`-.�8Jc��ke���n�Q��J)�Z����j���8����������ϰ���#�C~��ޯEb?�g�M��6W�Fx	�H0�)���s�(�
���w�N��)�_|ui��j�����P�Yi�U,��[7��\v^�O��ALA��W"::]��6����<�d�z/f���E�MM���/#���Q~�+ �mK]}])�����1�����0	��p�FS�6L��5�����!�N}�ԃ3�(Vn�$��
ނ4
yOe��8�\k(�jٝpAu���gY��}E�� r{�g?�w::�: 3��[3�u����Hɾb��|Ey�Gܩ:�s >�4�~)�vV����n�~w_���>��20;Ȍ%R��M#C����y2Fd0�l�[�M����%��Mܢ:���Խ�r���gr��`ԅO��W=��e�'�!�����8��ag3P&����O�?)�^ʂ�����4��Q�����HXǊ�3���~b֒�q�i�j�R�FSA3gc)��}��FO��������dۭ��7D��p+�W���#��S����)lJ>�L��ؒ"V��Elu���`�*5�:I��F�ǱRŒ��{@�����&e�!�$���J��o�q*�8�s��(%#G�=�/gb&�<s�����ةR��޼��T��a�5b���<��_훑=^��r�3,m��b7 vV��i/��blV����/E��AR��O{�F�Tx4���^�5�٨����?��=8]�x{N�BL��TٶA^��ˡTY�)iJ��Q01�]���z��K3jY��Mb�F]��ll�-�h55�G��PiR�Rj]�Z�(pf-���^�=l"2�E��;*fw��w��"E������G�yA��=��{T^�ϻ��N�t�w�>#A�ф�BN�C�nz�«вpb$��S�A�����z�l��T�����#ˀ)&���Y&��m�)}Y�H�h��(ۡ�Jˮ�W�l<ZuN%ͨ[/�n����  �#Q����:5�/�c1.֌�}��%�)��v_��]��Q�m{!�5��;��<a���X&N��p%#���WCy�p.u������Ѐ�*����3-Ӟ���x�.l�#����)]o��S��0W�dR{4F
U��Ѥ]Y�5����$��>{=w����`[?uc�'u�FE��uZ;n�.�'���� �z��:�B�L��U�o*2j�!3�����oԩ).�3'%b�)hSÿy���1�M�%xwL��gz�*L��"D�Cl�灍7��2e�h��p��z�/�i���h��3�Zޖ��m��TG�[�?�H�n-P�P�)�r�SU��Ը�bJ}�ܬz�j���[g� ee�~������;��Z��,N��� ^�C����%�������ݜ��߁�'�mx�_R������ϵ�Ĉqw��L�:�.��
	�5�2�GO
X�vd�1�~	~)j>��|E9����m3Q��Xޞ^������'ĮHh������h�m�?�?�!�wn�	������*�o�w*�[�8l��y��B!!��l^}G���ZB��Ԑ����X�B5rޯA�Nk���K݌�<(��e����8*����&�%V�7��]���.-X|�_6:���L�ZU:�����Z��)�h_Ș�s��(���I����zxu��u�C_[M9���{�Yi^6ٿ�&lH�qM��$9&'�n��2����0|�aA��D�7C�@ϗ[�)<�ݣ�2���چI��$1�_H�:�b0D7��5bN��1:���?M�>N�s0d�L�ŀt�ش�z^]�Tx6ϋ���q$��QJKK��,�Ԍ�؋(_�@����d�&X�������+�`�z���j����LI���q�{�G�'%���T�ˆ^֧ړ�u�
W��x(uh%<9��?/>���i��O�8h��GxJ����pD�Ö�䄒x��W�d�%�U�JA����5�[Z�OM��� n �?]��7\�[�}�$�x�:}�%���:����3ZN|�&?Y�Gt@^�Egу���Ku������V+(�	,��E�lshx��q4�z�9�&ͦ���֥˕���Q�yA�I%�;Ct)��
��Љt�g+c�G7�CH�7�����5��EC��F�h���}f��������s���wF����S�Y�>G����f�z�i�!�M���l,��w�h��+�4oMY�L����y<�����..�l�c
*�������@Ǖ�M�}��O���sЂ�
+w��U ��
�J�	q��������u-�-7����pp�4�	zN�0�I���c_;?���HJl�rK$�w0�����b����t�t0`j-l��A��[l!��=8 �J2h[�lsM`h�;mY�v���R}w�i�� +��4��Ҳ�a��n�>W:(۱il�P}j�[����5@���2\DN�qU��? $y�7�S��q�Y=��X���E(͞�8VD+v�,0��D;x��m������1��{���1Z�eEGJ-�h�ka�kt��+�ߙ/����s�ӛ�U��
��T�&`����yLd��4U�:�E�sVʩTQ�(]�B��[�/�7� 3.�i|�8�_~$48�ǎ/y?߾}�8v�?���D���F����x�X>���<nV��zD�I��wh[��x��pE��lS�`�j�H�)�x���M�`��n4j���M:�Z��L��RHΊ�(��Y�9fўc��T5��R��"�t��fh�1��`<-dJ�U`E�z�Z;>��d�]�� �^�9g~F(�;���nL�9�ן�xp8/U���@A��`Ě��P)��@Fi����"A=z���Kg����`�K�ab�[{����12Yހ8�$�n_�1�B1)�.<کk��=�JW�~Sǫ���y�bJfpȉ���� ���ZHJ�,���9L��Đ���S�[�C�5+U,X�.��"88jvU�����*�lz��������j��(�|�a�9�}4Po\�M�g�(.=�29Àí���cl+�M5k���ג��Ŷ̀�-wy�ޕB�	��%���)0�R��Ba3��h�Ñţ��%ɱٗ�m�g:|�ǐ��D4���ZS�z��/>��m�M0�b�-�u
�{*���	Z6V�WI`�W���]��8�OG+{X܀��A3K��p6�㸮�P`>��[��y�.ϥ��׽OF%�)�}� �\�w����[L�w��z�7g��Ae)�=b��4=<pe-NpQA���t�j���;^��R�=���f(<��#�ō2�ӗ�<R|�	�j=�\������(~�2�tO6��Ϻ�aO�"A��Z?)�����ɸ)�O1f�B�2�Ԣ���P�#n���� |�`1zD����i�;�Ps!�h�p�M���"�o����$�� 8k���r��8P$:z�GYS�J�6�j��Sy�D#¡TZ���~D��m���Gk�ޔk:���lǑ*ׂ0!SjP��&m�^I4��d$�1f�e���Fҫ	 ͖�6�ɥQjV�Y%b�%���`.9�t��,r	�����J�u�fA?=�Տ�Y��H���9�%�n9��Jv ��6	����5 $V�7ځֵ�UӇgI	~f�|f��^�X���>t��v������
��R�S�eI�^K��lnW�;�Ć�[��D�@��>'��eYN)��%���<*��}Ywj}��|�`H���Pٿ��Y��V<Vh�1[���Q%�b25��(+p=Ct�Z�9Dz�{�����,�/ͭ��S#\N�犎�ev��
P��hjj�sʡ�,@����7�a�+�Ի������l	}
���T��Q���^����:���=d�{4l������/=s(�u�*�I��m[�F|T-�"~�̊a-�,Bt���W�U�eB�l���W~h$��:ɵ}�M�����U���9!�(pΣK���^�_�7o:)嗾϶��b��h��=��Y-jo�!��'rdd���ͬ��a�h}G���b0c+Ɣ����vD$b��8CqC����Q���V��|�������I�%�� >u1!��d;j���O�I�4�p�xi���({re���y]����P�'j٤�=�s]";�����>��嬳R����p�K\V�\�������6�'����Yw��h�B���D4ky�q{_��rF�U����d��˟2=V"�Al~�Mn1)�돔H�� �l��*���HL?�vkqM*�=�@���f�{�;���ǃ�G�~/A�.��m�%�� �"�w���%cE- ���rg[f"*5�:���lm��}C�V_X��L��ͅm��PE�g�	zҘ��v~�^�X ��V��#��8�e���;�Y2s�E>��"��k�����J�P����{U��g��%�9S/S�*vX���[���V�Ü����@��ѹY���\-Κdg��VN_(M�_k����[�&Lxf9��=���>l0p�A�,mm0��ЃiA�f(69���_�X���-ɠ�O�^���/�!lS�yP�ʏ��;Ώ1bV�Ց����:��}�J���!�ӲJ%���	�sE��k-`6 �<�u�wZP/k7q-�)v����M�K�˲77��J�0ů:Ϥ��G:��LAjN\�9#������e��,��e�u8��N�㕂��R��G]z0+S�ܤ�v�Xuw�ኟ���jLn5D8&�S-��X7��M�TD���:A���fZw*��,�S�p�ЧX9����s�lj/��~����N#xOM���c��HwI�jdn�J�o�:�9�K&�o��T b�.Q�f�?�ؙP�ke R�3�]��x&�P�����ߝ�l�sz�F��U��2�tU��E�U[���1��zA+��TKO��$�F�p	H�P���!��E���׹�3H�Q����C���`C���֨�I�H#P��	���Q���+��t}�j�e��!l�$L ��xXw�p+��aj�kb��s�����`g�j��6B'�5�V��^��	K>�"�sгf�{V�J"DDaO���$��=l�V;���6FJ�5)3�c'�>g��~�~�r-*����R�B�3#䑅0[���`��]L��8�c����FXj!`�
�3� ��,r�\k9Q�N2�μ}���Hb��C
�E��l;�΀Ɍ7$0Y8��!uBXӾ��G+b��':z��~L%7�Ʉ������[�B�L]����J���"�}ۉ�j�\ԛ��@��p��N,?����J�G��c1��T���������l0�l��kVT��enS���������"Ǚ��a���X��wFr�~LB0��E�/����E� �\v��\Yzڴ�*�QE�b�L|��痦������anW?� ���:��!�;J���em�췹�Ы��(k������;(ߪb��v��K������Ĵ�:"�VUޑ��@���ᚰ��I��-x�e-I��}��y���ƊC��+p�x&�Pe�{�"n�X|�i=�`sG�<��D}c�vMj����F��<��7N��a�>�����o��]�Ȧ�?6�飴/3br�t0���Q�A�#����ekd��l&�	i<E��4#<v�g��Ip�A.�IK�{*����Q<�{Y��φla�Q��E���!M6�j�����c1a�fi�<�W��Ev8���� +��jVk�\E`�ʮ��Ĵ���5�z�GHy�,!J�����Ú�N��z�����7��ͥ��V���Q�Jc��BC {�d$3�::�$�Ǆ�9S�@�w;	`�p��qD���gz�ʤ�6��ɏ��ǂ����;�b1���բ{-�ش�[0�O��xk�Z���-�#��BW($��~�&�+��]�[u=��d*��l-�7~ݕ��ٕ\N>�q+�YxS�O��ж��a�.���_���ѱ�/���^��Z�]�D	 �㯴�ѩ}]�t���{��vQ�M�Hr@�'�f��m�� I�o /t:����>�<�ʫ:�G�K�Q���g�/���̙�Q�+:���OҨ䋷߇&�����
�Vn�M��;�����g������R�I[&�����D�X��K���	
�דXY�L�l�	�/n�l����*S����ڰ��������#p��1YD+��{Rrq���YD���2��Ϊ_�u���d�F�h���t���aU�:I��z�y�{����P{K�M�܍��)�F᪯�|�C�����W%���7_kt�=w)Q�SM�K/�������Y��>����8b|PI�w{eMv�:���_C뤑�JU��n%t�_�jMQ2U	�F��g��iȎ	g�:��K9�,���)�k��w�U��Z�tm���'uB��3�r�L�o=©ڇ0�e��Q��*!s3ky�ч���.Qur�s������F=������bZ��٣��%�|ܪg�J�s�����D
��kW-��s�A�X��~�5W4z�2�pB��G=��<��J��{�!��L5�í8���6����w��W�m�j�ܲN��;��u��;����N��[�N���_��FL[]6�Y�N�}cu�K�_�� �A�-u�N��	��[�c�|'�t�XU9��@58�D�ȭR�ŭb����X;6ug"��Ļ�_�������#fM��t+X�!0;�r�C�Z�t�&_T�T�:��9�-�	M��^�`�iP�Ɍ�_6f C��5М���9wZ�Ё� �:Ȭ���w_0/�il#����$�L&����/{�,f�ūX�$�ҏr�J��K_�3-�k��N����O�KxD&�}�@b��<�Xt&�;X0/b�C���4���X��C]���U&��?����y]�ٙ��<�@�>4\88�4�(���%?7��z�'��~��>���ݍ��)WE�kK�F\Fih�x_�^'2���ύ~hm�y�d4���$;�I� ����g�m���.\����V����#���߂�E�&��]�9��{�������٨��z0���ń��.+��C�����J�譀9w<�