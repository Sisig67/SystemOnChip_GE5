��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���!<So���2��E�!�7���feI�R�34�F�\1uR�XO.P㤳��"����(W�����Y�us�'�V6g{���/�Y�^( ���Ne�[�����8�1��{SZ�k�eZɇ�FUHn�i!�kO����r�o�40e�@�̺Na|�g|�O̲s����_�oW�h+c�	��x�1C5�]�`��P�#�Ι��;<��C������^c�4�\us	���S���x�~T-���]D�lK�c/[G(+ف���j�H�3!`��|�V�k�)j���Rrj������+!�m�iS�\�,�D nP>�:V0�(�9��O�Y����m���7Ӧ�J�Ā7��-�o�6���d��iP�2I��5����^��1֐쬳پLƑB?�(�x����wj�j[p��ب�Q��8�)���b' �{b����Z�مIt<8�3�\;++�Ҭ���7���$5�?��Hf���*"��6u�Ea1�Q�g=�f	����%'(�l6���g�L�YG9�:x}�� ?d,2+5���1;T��U��Kڐ՛vN��~ō능���d�>��$�s�D�Kb��{��V�L����+��6pM�ld���v�0f3���w�ہ�V����W��� TB�Ov�4T��9k�m����Ҟ[Cṕ�Q,:/I�ff7M�d�$#*�=չ/Ȋ?@O����-�+�g`��0�E�΢f�Ր�#��l9LBi�-�.�{��޼W��������Jx�a�8T�r���ŲG��@�.�f!`¾F��^~�G|�v �FLN�j#!Mʤi��ɘ��R�������L�"��[�V:�(V�R�Н7�i&O��Q3��������>ac-k�cq�"B3Вa���-D��+�;�IYd�xޱ�T��F�A��Ji	���π�[�>pE�����ðh7�A�P5�f7������:��_m��\󔊁��?<���5|���b�P$1u� �,�U�����Q�	$��/s�QC��Tb�����nO���n�E.�|�@��}�"�^_"~B��F͵�U
�Zյ'��^L18ik?p�:�yo�K���&Q�V��b�՞�	�Ja�2��ň3�����c�R����k���+�T���0\daQ�E��B��󈄃���.��mUו�h������H]Zl��+�"�?����hK�;�URY���v2��S����y!�	ѷ��7D [���~��[�?:�����&����RT�Bo4)�~�UU�P���j̆�j��F�4ёN/Z���q��8'u:�|O��йIJ�f�}�":����Ep}\35)���W��.2_�{֔*�~��U��Ȏٻs��9���ɍ/Rl�6T}�8����
�%cǫD�1 M&��9+��^Јa�lXoؓ�%��S�*͕�`ZH0�+�D����;,�g���m׍~�'�����\�E2�[k*�,��=]�j�,w�u!%��:����{b @�Z������t;PL��W_R�}�����9�����T�i�z�o#	�=�
�K|��<vx��;qe䊵:&
j�)+=��!��1w�G���yA;�U�9�h?��\��L����^��gjO�Z�������/h#b.�T��J��홱BՔ���Y��UB�����)2.@�����zb>3��J�xӉ�K�c�aNo�9�@g1��X ۇvԧ���2�W��Q𵛉�5۟�K@W��B��tѬ�8LH�q��os�� 0]�c�	���H�?��*���H� �͌U�D�^�tf��n��@�Z���U�IY��%���*�� Jt3�Eүf=�y��`�j�s5��A���W�N�?��]&��4�N�,,0ڷ�<��kp06��k�&��C�?�x��üG�^</�F6xw��9u4���US��Qcv���ҹ�e��X�W{=`̴�s'L�״\��{D'%�z4�E��� �0�Z���5�Igv/�bn� 1t�n|5�d�yqA�d~��p��5��{4*�_$�Ax���O�ݑuI~��O-o�A�-��di�+��.^.�����q�6��	��l���Ə�Uo�)b��ft���:��:L��`r�� ,��ᡋ}���4�w6��*���G)Nٝ�6�y2�4vQ�ӘT���]�m3�f<@N-.(��}[��=> -+Ϛ��N�i��଴A(�W��:�&���X�}t��U=!`G�A]��Ⱥrl��5��)#�38.��B��m�d������*M+��CT��h�;��Q����s����8*���.r������?y3������@?
���^�й.ie"�8ü��� �U�x#p�@�����W% ʯ�ڏ�Ti]�ߥ�L��-��e"��&��B��� [$i���kG�����1���3; ��ޓ5� ��Ջ��~_��2~�VI���A�:x�o���b,V�Q�����D=�'&��%�I���`҆��uQ��hh���˳'�	k��Z�\(�B��`{�.��!�ц�
�?�Q�n���00�Q7�:I�L���N>s!E�P������.G����3<V��=���r@a��u��E�h�Rq4h�o_���1F$v�'F��*V�+��5��52��y)��L��gLĎ��,z�\�h����=�Ͱ���P�ԡV��|��~,�si}�;�GBo�1�g[���Gd	rQ�\����EAKc��gks�2�	�-�J%����K�S��EfZ����q<w-5��8�()V>�%�n>�ķ����En��z������0���$��2&�ɸ�C{�`3x�������YY^�X3�����ix}�پ������w�6^��^��0��"�e�wxg�����%%o�B��N9���Ҍ*�>BXI{���	Ђ������lx:�`�&�r���a���x���EH�/96o.m��O�`d?	�j�ZWs�Y�Ȋ{�N�mbb��k(:�C�Ga��VH�h��nZ�d`��K��4�� ��u��&#[3o[sUkrs����a�����YA�B��zx8�h�c������8�E �y������pE�
埅��O�"�����ʝ2x���o��D���^!'�C��_o�A�4A�%>��|r@D�L�<���m���9��-�D4�`��׿Xr�Ɇ�nc���^�����%ݬ�S���KBK�h~	j�_��.q>a�V��ɜ}�rb�S\�E�w R��|e�xv�A������xc��taS�)�E{�����y�6!��=��� �L� v9��:�P���Y�vuFB�X���v�[yc��c �y7�௰�0�J��}�M���%�E�2��j����1p(K��+D�}t��Ō�>�\
h a�Y`KP���|���o�"\�_)ʳw�0<w��Z6gU��V�e �Q�(B�6I�6M C���吠���m�fB����j��Y뫸*h��#��
X x��#f�Rz�>)~�S'�����r��V�*Y6��a�\����8��{]��5��E��o$%�;����=\�:wx\�B���+��.1G4�}qҶv]�u��=�ǵ��WW��Uc�2X�:>����^Z=6
���%�E�9�*1�:*�=e���Da�BX�]�t����B̝��b���(��-R)��i���Y��	�D��"�p� ��	7|�
}g�#��T������%i��}���=�P�D��w���`�<�SG'^�_#Μ˹��`�_b��wY�?��Y�IN��`�I��R�������[ȹ�-�\�0��G�2�met�x}U'J��Lrᇪ4t�kn��f��[y�P�7�vv� xX��v��SN�_��bj�J��6�����*'�$�g�/��y�i#��J��)�'����A"����	c���qBUǪ)��&&%q�?�j�9p�����o��ʅ_�a<��ִ����T���B^#A��r�b�yi��XF�����T2ZE�T�>�L)O���}��r���|�tv�Y�%�9g�ѫJ���=Y�Z'�ˍl�X�ˏ��+r-�P�I���w��ǻ\^y�4���e�y��J-ᶑ��)Йo����n,��0n���Cz��k�2��LnH�J�'BH����L �OE_��x5���;���U
�gY"��	����^��^%����0�h��E����N̯� QC7���Gۚ��\��1� ���% y�h����ާ3pUկK�
�!���RP.>�Q
m`>
T$�tG�2���S��L��:�
d����7����bZ��\����^�?�bѓ��hZ���(�p6D>��yc򖄶�ӆE��aR^l�SO���j����g�����czG�ӷ�U��X�T����
�L.H�րN�����C�i�`^�t��������3@q�v�޽�\�G�BF���1� ��[1��C�hj7ab`����`�m��xA �Ծ���~��b��|[��.㇘��r��H8����Q����}����!9̓�u�[�H�[�P6�C��I-��	L�����%�,���-B�V
��\�b�o���I��E1�=}�� ���@&.�� �D�R*V�tJ��)��${�V7�<��_�����t��<�|�ao^bMi�~&�͙hV^��E���t��(9�?和X���D"����S�����$[��B�z>{�Z���iߐ9�x��ͬ�V� 0st!�����0�ö^I�Y� ��sB!����	��#���5?���rb�� ���MG����r��?�ӟxR���d����1��o]t�s�9��;�R����nr',�O�?��S��x/=&o!��׃_0�b�&��}61=����e؞���ɛ(����	P�bt<�#vӹ��oR��'�[��N���p����*dysϴ�6N��Ѥ����<>y�R��t�/e��,���|��>�ht��u.��w��^��e �S���j/��2�_D{��oJ�ܢ�=�?���/��k���uS�)�=׋�J�Z�%q�@��g!̪�sR�_�ƔG��Z�GҮX���mm�X����?ۉ��Zj�>�?|s���n?9~�6 &��_Ep�� \!b����4��*�R�]D�3�.V�ׂ�>y����q�F��x�n�I�.���8^(ZI��LQh����ҖbJN_�5�S+�mBǈ@.� ����z̍�o�2R��~qi�&��0K�LY}m�����c���;1�Y����ĩ�^�V��.u���JCȶwR�5�Q_}N�{�ݭB��y)�=P�?C���qN@	�E|��IJ���,�_�ذ���ns�P�8_�6קt�*��B5_�~>�?l��:R���j8`��e�ڹ�(���-'P?��U�s� 0��۫Qpa���g���r��z���V%0G���Qzd#Tc���'g"�R��;�Ӯ�1U��m�t�v��(��`e=C $��{S8v%�*�H�XL�.� j�Z�F���FG���G���!�.�,����9?�k��>r���B~� q�!Һ�."E��^zX{Qoj���.p���;��?���ܮ���5ʑ[��Iw�Ѓ�Ͻ-M2x��w�`~V����gx)=��\Rt��~ԁ>c��~�!
�޵����ZX�Fb+~�#��c#Y"5�*!��$�E��+)�{�����ʑ=va�J)Հ 40�G�� Ѓ#n�6!)�!���;vN]�7t��;��L־_�N�
D�o������CQ�6�4O֔*��S<
_��O_��\��fIb�}�y�k����ց��;.�+�.1o��s�Y�b�מ{�F�W�^���(�%�設�֒��J4縝�(�+� �	��-��6�YO�2J��}L䐭Q�'T���m�s�^U�N�<��\Y�!�qq~b?|a�⃥p���ߜe��9ݶ,�M��[%�<1�/#��|�x,��TLҋ{�jKI��[� od����+�A>V.�zO�O�̇��gBR��Y-f#N����wG�H�����[Lh�z`9�M�h�7x3Z�1�ƒY8��я��
�������_��O�=�(g <T%���31ڿ��b�9dS���
��!���8^����aJ}8(��:%z����y�?>���� 1�7�kX�*tIᨣܢ��-F��z�t�3�t�ﴷ����T�����[3nK*ɤC��V�s�;�mr���wB&i�Ux�m~�R����8�kʠi��ƛy#=bb�����o}����i��An�c-�����	گwl0\|�h*h�H����0fE ��?����D�;�z����q�,����pŻ� �n�`٣�	pT��[�N��p3
6��{�'D�&&�������k��V	��z(�,-_�<U�|����\3d+�� ��3D:CmCj{r?��{��ǭ~̎�g��b���F��xԕ��k�3��M�'����!�ʱ2%�>_rY�oy�ߡ`�m����?\j���V���:B��9쪊=��ICc1&��y
w������I�_� :�g�iF
d���-�g�n���%zs%�����ye��:ʎ^'�8���Qe��t�;�����?���^f�/9����I�=��Tsl"��� �d����4��F�3�A����b����SS��M��)�����^��
�����S@��MP�#|1ũ9��.�x���4��@��ūx�m�S�_5=�^�Y���B=�&�4��:d�O^z�ɡ�� ��(�߭�]�,�����l�1<�(Kx��*��9Xc��3K�E斮�M1�BF/�#�[���
�
�NE:)M������ۛ/�v/|��`��G�����T��u
�W���'���k�*�6�������X�U�!��ʐJ>>���M��B�ʂn��:Kl���q�T��
cX�e�H�����f�Hw�sH�)�*�Wh.i�M�9B(��!��UmUlZ-ٕF#X�s��U��#=&td�mQ*�+�\׮���h��$�����n�*��청SN�N�HGP�뎆zW�FS�Zij����d�{�Z�G���P����/��뱱���˭�����u�5�wB�Gt�.M�ԕ*g^u.�>{�c���X(�~��J�n_ί*��m@ՂLBUHh7u����g��B�Yt�������`nBE��\흒�&��H��0S*~��F7��0�Z�"�Co�%�$*��gl2ۏ��d6��a��+(��W"i�6v�n|�ZGk|�\ ���p��)ބ�'-��&3d��kv0�n���}����O�!��'�����[�i%F.T�q�ȝ����?Ew$�.�!?�C�UtÓ s�e���� [7��>��un�xU� +����p�kh�����f\"N���#����������Q&K|z擸�'�;K�\טKp�l�Kgbqt�қ@g�x}㡗�[��n5�UG��ʗa,��?b�B�(�;�e�j�r��
Q�L�+t6~�����eu���4E�՞�$���!6�td�d?K�y�z�2~=�5�]�N���ￇ������~�l�R鏸�c(e��/:�k��� ��=E�!�1y�l3��0���Cӧ�mrS�7�c���=z�,����KB�Md�a&��IA�]�u�A��:&���� �I�(����%�%l��JƮ��,��Jh�n=n{�FY��j�8e'8��O������y���!n��\��B�/��,�Y��a+�I�%��9�
�	LxECp�+��W�h��2>/�cc��b�}�*J���~���P�L�i�L]�$)\�9?�
��k�/���=̆��Hq�]��7�o����n*���7g3Z�"?;���M��	PHO|���c1�A�N�E_�[dI#� ��7Q��-��@m��_%'�P�4����[nJG��Ɖ�ѷH�ł�y'_��K��17���3��Fcba��ӷ^N!�S#VL!��;��ޕ����y��S>�VK��)���3�gN@%	x���,��8�	ѣUE����ST���/M�)�ɡ꾊�v<�D�J�g߁b{��"c�Z��:]*���<໬���F��>���{��p�&�R4zu��k��߂.'v��g3�<���Rj�߄V�FH���������@���nv�n���$2`c�;�|WHc�]�[�r�ا�U0֬ئ��;ڞ��Z59;@�.̚H��|����ȏ$�N	�pg:.�d[K. '�s�&��nv8Q��74�P�_��a<�b,�l��\:��������E�u}v���w����`�xߞ�����w��?(��tA���(0���	���?T�r(��ڋ�P,y,s�
��	v�S�|²�oTf=@?������*�)�e^	>��<�A���S��1�2����)��eՙ��*��S��9\oq�h�%*���T/[���:e�sx��)�����
�Dx(dG�]IP'H��˿�g���՚���O �i��޾��vf�Dg���/�׾���n_��]E0C�mVO�sIg����	��]l b�bm�A��*C�<�"�J�;��a�}鎞���l[��<��B՟�X��	�����p^�pҭB�q~���WZ�%*�RN���s��Y A�ӷ�r�{9���!��YF�J���eUI"$�ڬ�y6�a��H/��^Y�ب�tɹ9KH-�ڵ[����A��E!�+s���9���d��E�;�'�n�?�E��%��E\���k��c��*`n����cE����n�xQ�����G��5r�.d��Wg��'4�!�x��,��EN��Җ�8�#$XQ���E�V�aߜ��RO���Ιx�HS�iM�Ъn�z���QƜ�2��@���4g�`Fp;zH0T�  ��I @؍��͋ԇ�#�����Y���q���z�؋Je����6���b:�L���"�����爕n�m7swF��y�;�H�����HfW �9�a�W�~p��@:��*���g-�
TUp�ز���)��FړY-�q�V!�4p���?�$6��φJ�x���Q[P��KJ4/���ۚ���#��&�N_)����z���'�T#ܣ�F��E�N�z�����u>d��)*ekۉ(�k5/�m͵̫��$M�"�)���Ǻ�M�_(/[7�7o�-\�Hg�ZU'���`��*����z\�ʂ�P���=��R׫��XO��q����fs�L���R.]�y���㩱���3��ޟ6�d��L#+�����$7���1rql?<���d�Ԡ�k��g�����}T�I^�\�z͡b����VI>[b�y�5�T3ςv�I���STc��ݞ�!��e���
�r��M�~$��3�����JŞ ``�mawhi}0j��o�/Z��b�G���;Eg"@�n��3`<1]b��sq�fgw"�YW�DtX廡��Gr[Q��F ��^Da�K+2>Rܥrd�a�r��󶇥k�q|I��tQ�0��xq��)���s��x���gxy�+�F�<�M �U?cd�k�k�ֻ�.D�~y<#��5{�>�Hΐ������cC��E�[y�qU����>��
�a=��:���O�C�����3u[�3@~4��x�&2ǜ��q��_�������1Mtu�O�1�ۀ�Ōs#y��l�(|Hm��HC%$\й��0$M���"�To����}�g]���3p��Q;`5�z����4�6�p����*xh�u�@w���N1h� �� %v�LcuUS0�����D�h|�&E�d�S����֚(�!��fAs��r@��Ds	Âe�C|�oJ�s^�k:+�Q�LU��;?N�{V{�3��Yd{��ΕhN�+(�S��*�/��T�^�wA�~�\����+y��i�aެ	`�ak��A8(rE�,���!���JIB��:x�V��l3�FYw��y]_+�b�NӨ��7�|�C���9��U�ӵ3�=����;m��d*
6�u�KӇrQܦ�G$M~���3P���F��=A�3rl�AX��4n�2���~���,j����s1�Pmс^b��sY���G�*{���{Oj���Y��1��D��7��\�z&�w�lGc��� �GG<O9�YE��]410�e�1J��2�|�|�N����G����@�Ya��*�2�Y�o�(x�! /�[��F���X�^�݆�?h��bM�M��88;�cJ�H�w��c$zpo���S��]��J�KŶ�<��I���n�H딾��]�q����G��'1��4�
o��l'��}�i�+7N����<,y�9�,�z�*�|���{d� r�Y��q{�-��Ǫ�9�]��� #�F�o0)��ֶ�K�u�;�W��ó0�L�bç{i��ú@�Z�>���N#�/��3���V�i��-�Zl7㏊���:�sf �f���J�(��'��-�!;S�9��j鯂�M��"�G��!k%���i��t4�N�|3�L]��לkI��G��ֱ���Ә%��^[�Ւ"K�]z�B�W���w��I7��K<�>>ͬzkm�n伸��7��c�6��F�!<w� F]��j�)�b��DDv�.��Y�H�m�5g'R��߹FQ3~����$i�P��b^�f
��y|�Y���2o�y���`(Yř��u[�sz�]�M/��w��Q6���%LE=س��5رdV�t2$�6u�gw`��$bI�'��3�|8��	���K�I�4��(ԍr�s^���P{d͙��*��p����;���D�="Ge��6tj�DzlXmxp���2?0|!�O�cRƫ�GKW��o͛잁���^	��Q�%�X.Wr�PskQ���]�����[�G��&�� ��Uj��������[m�������KK~���)�q�I�>�=�C>I�%:�Yd�Ý��k�<RI�ݽ�˖$1�ؙOnҀ2H�1���(��T,N�>�-_�A��l/�
j �9"m�ޓ�ԡ��t��{���<��W]t:{PR�5��W1�c���ЭF�!HM�����ؽ��Ѳ���'C=+���f/�D�2�\���=������9��rh�-�#	3������a|�U�dj����zX���'�f6K����U���?���P,�N�O	����7��;��T���l6`jJ4�5(�h���w+���#*�ugʑ̜~'�×y������ެՙ��X���r oWo!mit��J���i8�Vb�s�L-Ќ9�c3�M�i܂��L��lh2��{�y4�X��,�eg��@#��R���;m���ޒ�m��	p�o��
6����d�k�-vB9���v�ɵW����b���j�.1^"�4�vq�l���9*��:�LAQ�� f�v
�sM�_�������_U��G5�&�����ѻS�Z��#̌ȑ����q=�+�Y��-�H"��H��8�iV�z�`.$8�M#7�e��T2؋!2���h�|2�3����h�/�KVb����2T�d�k�|w_<1 �8�kz@�.�?W5�F+�n̒]֟��cɒ���9��B��C�R-#�@�/H�
I謍�� [f�!#��c���C0'����X�ȿ�����<?%Ҭ��� _PR(]κߗ%c�`���k^p�SO�u�htq?�_<��!W�:��qw��TZ�O'j�z�q��?zg���]qWcw˨�bǝ�oJ�t���L�u���(��?q!(�[��M�
�5����������j�����+	��m��7x@%Z�f���l	1@�k��;ը�ڨv*; ���!��zKO�B0�̈k�;e��#����6��8�_8m)CU�~�%�Uɤ��g���e���.�
۬�����a�o6M�j����9�&��$wR����r�Yl��%��w*�H[Vg'���%Z��t���g�t�X���gs��.c��`�J9�ю�-!
g�)�1����ou�C���Er��s����Q ��t�����`R���*�J5u���ɼ�o�v�F:�솅�U��JF����]��T�1�=у��*�[ֳ_Q����=��"�qn���[H|�e�m��(��6g�ƸY�$��kG�S�@e�G�%|�.�;�X���3�4y[�A/(%9�)&���H�\�5�����jZq��V�c��܆
�#[+���B rZp:-�v�ԃ&�	�&d��3:7U�:SI�gNCUp�
��c���19�Y��`�Q��y�04kV�-��F���6�I���Ut����S����@y�i��gR}3��$3�7!p�<3q�X+������,4��e�� 6����8��_&�I�O��ޅ�#2�W��Sk0gjí\��_��@�M�nyp�/p�� |�߼��$SA��<NH�P*�S��~��]�K����&�jT�f�������������V�bl�v�|�y�@k`�߃��a�w]�WcWd"�y�y�Ft
��2�)��% NV���9ic�G�α�H(�j�J��h�5¼��.����x����.0�͠�(j<�yI��C�A�`�U�A�o��������[��r>��E���`���`1*:B���=��i�-.޻�����ۅGŞ�b�T� �La�#̺��
E;ϟoM��$c��Mܽ�r��q�2�qZ}��9��vb�_U��8G�nq��D���JÏt̂z���Ģc���ʀ�WN�vE#���A鿇�QN�T*7�=4��I��m*�L;�G�a,0��>R���n�.�,h%v������0֮�׽{�����  �|�y*�j'�R��_��|��#}��d
ӣhE���z��ak�_�x���6��S��	�4�j\56�X@!��oRqc�L��~���;�
k6kp. D�$~��۔Y�`�}�P�/c\l�_��`6ɠ����t�����
w9#�pl �.��Gd��3��K���Q��bwu�J+���Y�Ә<�:m�S�s�q4���?��O�?SJ����8	^Ω����0]'�c��{��{�<v��\�X�B��{��9�1Q�T��P���IZ	TM�Z7�J!BA!gL���j�����l�0���yW۬��r&��Ǹ��,����3�0��l��7����s�PZ���zoIs'`A�^s�2���X��ˍSw�9�L��Hy9<�u��K! �ع�_��`M��?�[>��`ZěJ�L��"@�^��Ta��F�������ꯍGk���ے;4a��	�pf֒��T�����f��*��w�Ōa�v(�"�oB�"^#:$x���Ǝp��tu��X]}��@ �hgn
�8:��C��55�l-b���&�g�{r8y���D�t,�D��ȵ��
uE%����u��
���rRh}
I�-i8����$2ЛԠrG��|}��0=w������o��[C$�/���AK��r8�0r�Ο�r�����Vp��������5��km�~�G=�Z�9�:���^�����|�bD�O?O�l�ȿ��Ur�ʙ.QN	@^�w�M>���M�v��Gl��a�AD\#D[��ٴ�c���g�7X�m���(��E#���W� �#."����}';$da�*�c�Ԗ�>g�"T�lLھ}�+��0}��]0��r�
=u9�AK#�*�(1V���IIRJ�(�+��0�ϊ6�
h��d����;o�5-�����_%܉7��5���Z~a8]��iHRCd�>�DJ��R�`�9�Y�ݎ��c+���W�m7��.�zR��7��m�����n`���<ݓ��/����j���~�G�
p@���o���/�����>'E��1)w0<�v��j$r�h�XfH�@
�K:�rb	���\�O�Au&Z��h&�/[f���%�.]#��0�����3o�9پ:VO ��Z&�0d�$����>X�z�`#�����ϝ��b�j-�Q9�#������1� �x>΃���#��յhX]5>l�D�ik��Ld�q��Zu��2Kৢ�0�V�w?�g1��[�h6Q.*h|��՚U��h�Վ(!\���{&߹�֩�~�:B'��y���"�n��Q"��rXf�V���;�sx�
���LE��@���J�����A���s�a�X2��{�t.~�Ԍ�V�������wRGJފ(F�E�������Dnk;����t����\a����g6�o�ژ�<�9��M�����%%	:��ش+��v)���i�D��[�i�Jjp�-e�	�J�B��_Õ-����GZ�����u�$WR<Lb�	��f@l�e�4�rl�|Ί
x��9^��Z6�qoW�(�˵��s�^E`S�~̓�c�&�+?�g�%϶B��m��5�(�{�C�S���AJo}��%�s�I�7EC���hr����zx����'�\���i�U��M��B�@���ȁfic�|F�{ꈾ;c������D��:Ж�d���[�&�N~��Tٓ/��0��f�sǛ)�O�^�:���tI�YIb��"y陠�#jԟlq��E~��]��Jx<���`��:����s���
��c�ݢ�lA�TB�y��qD�ևԁ���_����Cmw��|�n�9�G%�R �Z�|	��B{1�k�̖Fo��s�C
�4��G}&Z�M�d�T�Q��Vmg�%�̟�=�q�:����tI����r��?X��hV���O�gJ��Ld�����0%�Y�t���O�ז֋ Tb/ "$���+Gf,�"j�T���N�`N%��~�9�F����r������n�/7�1o	o2"_�x���gi���k|�p�YCMU$���l�~���m ���-OV�p
nO��^��<^��;�y��s�?sk[�|�je�i��$����wG���R��%�'v^dN�������f&xF:K��;�P�l͊6h��� ���B�� ��O^� ���Oq�^�A��G��\J��0���vg�}��
E/��p
���M"�'(�D�%񜂯���7AL�b��2���s0z��Os�1�����Y�YtSH-ez��(븾�̢�9޳0������&�&I����;ƻy�^�R���;/�0�6K@�Q�'v�#U�P��wC/x���]OO�b_}&���$�4\�P�!�>�g��R��RPߡi�����YW�%�r��!�� �d)�vGv�z��g���U��蟈�OT%9i��g�sG-\��_Xg;��_Y����'�]�t0��p9s���p�K�� y]��q<o~�3C�4Δ�����[���z�� �K�I�V�}�W��Z鈽8����י2����h��K�u^�=�&�Z����ߣ�B)�h>��iF���\C=d.�d:@g�͓j�;�>K>2��xM��������|yd�E�5<%>��,����f���ר�(~!=9�$��}j�"|�T�#� !��X�B�(ܑF������_�@�@��=�3`��l͐��tWK8�!:L8�ҧB2�:l�4�q�i-`��ٵ9����H]Z~�K�����w�B�R���o�>������,�Ve��Y'\�'�{�"~�$�Զ����fqa�(vaN21/w�ޫ�����゘\��ac�E��j@�\ p�9L�����f4�P�u����փ��[R�:����)�X��O���6���� �
��~S&Uw�я|H���E��	}���<���(K=�Ey����u"tO
�y6&��� ��댸�)��yIL��
�D%�V3��q�!�+�~ <�9���2���_���@��j�j&D���~��/�6�����7��]i]��k��kx�X��C��ﱨ����Dz<>��"'lR�s.Y�뺙��W���H�X4;�H��3�+'U���X��?vf=S����0�tl2�䨘�s�V)b����������ư@^0u��`��Annl����/�ɬ�2M�$<�0��P�p3���5ʈ�o��Lx��;�����q����K���̹f�M�:�ڵ���;/$�+y�b��*��v@��H��9�0��V�84��ٸe�ޔ���m1����x@f"��}¿O;����rħ��%��i��i����OA�h��P �-��D.���}�&�I�y\}\*�ʬ�=-��aY)��G��͋,Z �<�3R]���C�2�`񨅥����6˒b4��ԺW_�ɁL�Єt��t~��E;���rK�Ti5і ��GPzy��j���7i��b���{(�"y��R�N���?JV����E���Y�z	�w>�~�
	d��A����~��<-��s� ������Z��X�为{�xz1��Bx�5���8�B��T�ߟg=dVF̯ �~)d�����Z92B�������sT8���~E�r���|�N�lBO>�y˜�����Xx�%jYc��Nabi��cf	�Զ��ܒC%>l*�_(���H���&�$���VX�6�%��V�9�O�'Y��M�*�@e��5l1t�ɤ��TQK��~+j�#ű~�k�i��I�`%�X{��oe�����\�ZK��	@�KU����[��rx��U�<='U��aͰP�~�0�X�\ g�0J�}X�Nld�i~�ITL~�_�U#bb�#C�S���a�v�����c�p}h֭$M����s\HOYs���|� W��[�e�q�7�P5��N�B<��	��M��aU��u�]C���}�����ؔȨ(*�*Mn��ʇL��*�/6����÷�=@�w��l�0j�%x���	,H>���os�8TryD@���sA���A�"\��F���$uH�>��� )��*�js�#�ܵ��J�RNk#��4�
��M�f<��@6?2�sR@�.6�s��5�K��AH�<s�W�#M�AA�Io�U>�4��c��!P�K�5\��T�[�s"��F^(h��5yLC>D~�l�R!�),�Q�y�)���H��r��F���W�D>��W�� �;��a��6��'��N�0�$�i�]��+���@�+"���J"��������8��}�wL�q�Fйٸ>�xs5�8n����t�O)~�gy�^ER�6m��2h M.��o��zM�-�	��|�X/?�_h穕���{z4�y�I$�<�=@��@�'�	��xU��� ��U__(�Z�6�>�_��.�}�Ÿ�DA̒�6~�m�9:�]$�yy!U�F�����i�+�aM�ze��.��� �_����L@����5�.�o���x�L_Dg�>���n�e��|�1��M��&����;dBԝ�ho1G��|	��|����,�. �̞=��x���zf�r�T�K�}G�� )����.�~t�ᢷ�G��'��
��ϐML���V���ł{Bv�l�ꈈ���ں�8_��䡕��e����E��g,�d�`����(2�R{�>F�Zbz�׿Gc��(R,�h�`�΂Uۭ����l��Fk�aWU���(N|�#�F?���֕�,'$
'�_-�9��9o2�
�#��-���󶐇c��Gn��C"�S� ��6v���-y���l�C��\�J�n|�������=�}�� ���Gx3��C���U٦���THᷢ&�����M*���"L#\����m	Ec��Z��$^��_<�9�I7m×s�R�D�NQo�pi)-��a�o"��\���? rTpX0���`���w�!m~��]�,��9�f�|�<�bj����,�$�s���4����_Ub!��F0�az֐t��r�W-`fC�H��+s/
h��X`��i���V#?�'�h��^~�ߜpAH�-��.���s����T���DRK�a72���E���G�}O�7���eK2\�2b;l_����?���L�v�?��;��HM���;A�3�Q9�����=�����W.�*S��1��A'6�pf����`�}g"��U�N.GH��S��bko�g���0��WNg�tXhh�Y��$FQ�xO����x:C@���Kψ�B3�jP܀��0,�p��6R"&�cTG�T���_��+Y�Da$�S畯	d(.��!2(����J���%ѧC8� M&�.V��*�	tU-4�y>���| N��'�KB5�a@DN�7g���X)%��f�AI.B�ʑ�8m2 {,|D������E�x_�M㓫��F!!�o��r������� �����L-�J�f�Pʫ�L\l���8r��FՑ[@�S���b|H�����F�����{%j�>��j�P����s��f�Pi�zX>�/Z�aU:ݸ������0�Tt��wl�_�u�Roի R\�N��Y7��d��W�Y[�By�s���=��ʥ�&߲Ҹ]1��}�k9	�{�<(��j�<��}|\�h��y���Dl�7��c�E��&�4�as�������| ��;⍛�u;Y<����:d��
E�!{�B!�:(Q��x��	�ި�/�_"��t��XT�'�
0A�2�����<��r��{��s�=;��
ʫxkU�4�9|�	CZ�*��÷/�����~/������� �Wu��z�EN��N9'��Y��Up�h���[⳻P@.�`$&���=z��畞�{H"�<���ao9������;�'(�dV4�� �����p�al�;��X���]��!�]���W�n�|��V�h`���:��p_���<�b��v���k��&']Ò�Ѳ[5�� ���Qz�3"Q�Z���g���,�|�&���}>�1O��Y�jB���3_3�5(Fu�$.�Ys���A�鎻S��j�L�����Vl�kӎQ���f��8��� �:7@4S�2�y��]��M}`LՌ��]nZ�0E")v+��%ߞ���L�'��f�m(22\�N��+|r)����@x�9s��%�*aHJJ���ޚ���;���C�!�e��gU���)�mf�o[��ڛ���~l������������V����̩����a�.��q�M-��7Q���$S��g�}M�H���D;�%0��qY�5���C"BO�n�s)yv����-��]m*����.��}�y)��]��T�Mts���s3.u۶��7�^4נ��6<<Ԏ"��c	�x�
�&�
]�Ol��*��.�څ��;���Or�r�\c�ʀ�q�e�a}	?#��<�/m)o�����.sj�6����)п&R5v9b��n �10nG"+�dR�G�d����$����BDS�_�"^��v�ON)�IU��^�f.��	����-H�K"��S	�=�n�/�_���V�[F��9�
����"u�
IB7_� Cg�1u���]Œ.ы$�"� 2��*���"m�zh��j�JG;����_"��w�_��ӊ���*u�^Ϙ��H�|�XBUƴ�v�v�y;O��w����чUؤ�l��I�4^����|r���ݩS�^*�ӈ+��k���{��ᦽ�g-����tnxY��<�a��xFl�TE25t�f��B?�<�6��5�g�����o�wbd�
&�(ˊ��o��#�^��;�QF����G�h��g�;���4w��@�a<^�O�K><�#?�
L�~���#��r�=��k��6�a��B\�
��������{��A�q�K�jto  �������md2F��Df����I��<k�ؘ��[OZ"g#��ץwے���S�د娬l���VO,�Ap$����զa�Q~����G#8�;\̺�,@��Sy��/�'�b�d�)q}�gni���Ѩ�~�Hw�q����.J�I�'� K�u�K�Nw��R�Etf�s�yDM�$8�T��x������O �;X32���_�S /E�;p�P�JY��h�Vw��`z�p�V��;NS�_8
@�f����B�O1%�VLs���V���n�b�F�(5�i7u���ښ �UdP�����,����W�����Fm_��GY�q�V
[�����UI�W�1����p^]�(	 M���� {�axc6�ԡ/�Cp��1k�\0�����QqC�-m4Xpn*$�f��9*�q�,��n�3[	CYQ��� x�sl�I��#I��H��c�-3�~�$���%dy���g���%����������;T���qK4OF����:Ҽ�����t�t��q��4���]D�����d�0��QS�_�l���2�7GJd/��Y�I�n�ј�.�b��{x�9��Ҝ� HpjpV8Ϗ�?�D�ۗ�Ǒ�S������󊸏�<��p�˙�?9�}H�Ž�u>.��|��8[U������A�� ���j�@����PB�A�4�-`}�V���d��IX���.���'�$"5��&{�u��'#7 �z5~k��W2�}�Q
�V���S~��:��K��_�q����P��_=Oޭ���y���]/�Qc��/�ҷ�+����Q7 f��t�������B��g]}Hdb�9�3v�s�#����q;��-��9�i�4��e$Ε+,�Zg|����v9�6k��fal���ǒ�(�Z�j�X��7r�6�Q�����):/�Vm,�{鯵�x�׃|tл��%��0sI�{be
����ۀ�B�JD`�����r���*�z&�o�9��C���PqǨ��.��&��_�������LHL�٫	ʛm,�7 ���	Yǲ5
�Э�6�n���3 �O��7!L�g��OEIAe�=X��_��*����&In�Dj|���#��|B�F�dĊx�"8�e�Ç��j�9gz:�Im�
{l1��?/u}|��g۬{V�"����������X�k�Y�Kx#}=2D`�7�sh�-p�f�����C����F��PX�� �U�0$�']"$��S�56:KM.���%��pĊ*�<�������޾v�	
���8dS}���qi�-�����ͮ�%�����9�z�\-�~����}��D�H��J�la;�הW�����Ό���Vn\Zψ"�d��̅#�����* �0��J}����jO�61�?DYfZ�E�H�\��Ab%��E^A9s�N�1:��h:=�z�J���[t|�H��!3)8���YR�S���;Ff�x��
�a����t.hsr�=�������wӽh��֝��c�
Eb���_�=F����$�K}ߋ䰧4�V�4/�.��f^λ����jO�.Y^v�8U����fP0�>ʤ�A�ٕ؁̉��N�%��<,�_l�VO��C�3{����#�N����r�����J�7�\�]a��}�PНM�}v�"�>�z�._/�����M�;mRvm�Wywi!�F-3HU�_���zI�Q�����	!M,55�o��L��� 4�t����	D/1J���㺙���2�\�_�[Z�^o�,�	ȴDsuh�a��s�}"��x����*���E_G����Du2x9�#K���n~�Zְ��M�����?peF	d�(9z���j��}�L�P�Z꫶�x��r���F�1���}�Su�=j�M�E
,U_9.8�t�s�@�cE�������CeAÚپ��IEX3p�K����� �
��2�����=MS�$f�d�S%�uN,16�,,�n؀}��������8t�K|���^�k�'>�l@!��)S�cIsa�����8D��Ƭ���O��؁Z��DJ�rRD݆�x�Q���6��P����L5���]	?�NQ��b ��R��n]'g������˕�c!�P�wT1�?���9�]����c�ֽݜ5��!$CK��T4��]8(�^*6�k7�FZ�UK�]9�_�˗�JU�B��矷��<��v���`��9��5Qи�c��[�]!@^�SW��Vq��b(���ր=�n�E��'���ah�%U
���[����V5t� ����U�Q�$Ѷcm��;�8����fzDnS}�p=�9��3��/�S9��%KA7%+�b��S�EV��fЦ5}�����z�U�(�C�&��X��!��\e�a����0>k,@����L��z��Q���*ܥ�%�5Ŗh���%t��E��(���zn��ڑl��7�3�8`�»�%�cZeK�@��bH�g��d~�{��a*��cX��0�S�
]����mN`vB�z�Y���̽5�����%�Y�*A�F1�՟���4#q���aP�#٥��.��t�y#3���3��``[�p&tu���=g*q2e>����3.��v��j�^�1��F��
-��r
����G��-���
¬n���d�����L�6IՔ�Fً�����1����ӷ����;M�R�Щ�h�	IvJ�����P�=�1�>����}����l��z����H�@�0���nbS4��A{�\�k�c�Rv�Q'�QX����d�\��9������cZ�YV����I�*թ���[\Z�����JT�+�Ca?�)�F~��E�D�bw ��Kg�k��>������%���ⷵ� �y��ɲ-`�m/1���NC�4ݛ�W�ہ���8� ;j�Ǳ�rA�1�a�ML,�<�b�-�{u�㘈����S�Tf���n�6!�	��b�^hs��*�T7��ȸ�x�7-X- �0X��v�kq���珢��������ŗʥ£�W'�rZq_�f��WX��JR,��� p�����3�e^�#;�	8����?#Z�[ N�ۭi[�.�e�k�e�D�E����~��ܠ� 2����������+Z��cY�l�TR��\}������)8~���4�t� �hd�"���d������LH��**D��Y}��z�i���[ݐ��E^O��CZ �F�T
��$�����Cɲ�h�	�-gЇrx�FUYT�,�}�s��%�2v޽[�A����"���uY��7��=��<P)?�r��W	�;s���.��m1K�u�~���h3`_��2lwN�N��3g�c���C-�(wL��MAd���IL������H�~���\*ڍ�t{��	{�Y�~�ފ���(�093�gOS>PW5�6daaŲwKH��ލ�@��nDI���7�}%�唎ї��8Y`��"�ylQ5r�G�.K؆��$�0%���B��f!�.zB���t+N���� ��MFT�R�vȔ+u$�P�W4�HswC�t7���ޙU�)��*��e�;:0a&{�3������{W>�"��}�8g��O����=��|�?㢫��#�a��Xk���'x��H�ȹ��L����%:6���;����X�T��b���1u�;�Ճ�)v��+���iP��NH�W��tf��1ܥ���F�����<pM09 ���6�h�.O�2j�3+W��!�jF��pߩ��rK�\-�A8�y}h4�$�<9ȓt���ZPY~]h�J�-���_�1��H�
�d��y�B�t`�L��yL9%�>:=�3�
:}jxj"~�4��=O�O �U��
7tFX�"�[����C���a��l<��w�J�%���Uyh�}�������RP��.��R���aִ��<TQ���cI�Z
��v�{��Dh���n�k�+�RÕ�F�3��#�`�92�����4�Ĉa�0y|k�аo�ꄲ�{��+�l.�#8�({�H7�bV�N�7N m���~���1�)+\&��^����ģ���F�8��懸�f��"���
aj$(��M��k�׍+fs�l0>��Q¡͚O���� �����֒�;M���Pc��/]�/;2WR)�j=<��im���X3Y�t%o#*���wp �w�E��\�֚m�O�H�`�0LJ��(���N�Ȃ��B��^���U#VOz����{����\�K�%F���0��+�`xM�N�}[�Ь:�`y�v"R��#��O�+R��)��q���~�^�%���������YQ��S��"��ds����31�sA�\
�6�XغH)�SKe[�$տ�f-��b�B����~R��I7?�������&23���J��]g�8&5�7D���Hj�i���f	=����`]�e�Fhe�k�i�p����V��+̌"�et�V�$�\a�ןy5H�d���{6���H�7n��k@y��q��
UKa����p��i����I/���ښ9����ʓ����B� ��er� 3,��"�7�&�K�"/����0 p(btī�V������{�x��_�XH�C�x�J�>@;b�%*+'5#��lE��o��9'������3y�F�G�E+ �^�X�-�tn*��tԤ:H�x5S��>�ֲ��B�Sr�y�|!�J��$h٤�^��xgsّ:��ܽB�IW�m+@RgI�6Kr���_g��U*�3\?}9�޺��+����fC�[2H��ᚬG:G cп+�-�ԳzU��fOe>�����ǡѐ%o�+5i��>�Y$�2%�ާ�����2 �M�z�Nih�{t~�������Wi�<Z1tB��7�Kߜ_e�vͳ�|)�Z٘�E�!Hl@��e���Cc+A�1��Ctl�]��VؑYN!���NprQ��؁�*�]�~�0͐��DEu���)n ��<��F¦L��U�Q� *L�
����X�v��c���=����1S�7_b�ޟ����_x�w�7:�sZ}ʛ�c�)oh�F�
�ٙ%qbp�,�bA���=V��F�ys�:i��ϒҢфԕA�_�ZX�R ��kZ�/���'�����+%F��]1�H B���K���ߴ�o��a`�!��T+'}DP�e`v�e�)Ώf)�Jt���s��H`k�M(�Ʈ
�,��kgt��NS^ W����sf������}�j��'����A�aG��IA�g2#����V�.���e0�/ז���.�ăIc�L�h���\�t�D/�s����k�/�������83��%�+�ز��r��b����Ls�h�r� .��g] �t�.Xi2�a�&�b4>D��S��]ق��_f̼u��x"��Η�UW9���
Z���1a4�+���J�+�{p�� ~*�@k`�ӺD��
fP���Tl���O˝	iX�<�����d��^���f�(�>2�A/0�}���¡�4��-{(���(E��M�t�j��2�Wӟ��<д2�ڡZL+�v���z'�Ǽ3~����J�V�	i�x��@*�� S��D_V�Z�~6}u�yC+�@��Z#�QKc�$�)���h����N�9�����w�Zۯ�: /vڄ3�S���X8�o��@���wj�/1)�8�y�h���7�a3?����an�2�����1<K,~���	v���E4L� o�Qkb_�
���������Q��Z�BÝnXK!��(�����K����<��R�@Ġ��й���
���o(��Pm�3��,��ҫ�s���8��n��K�73�_�'0��- �?h�'�3b�~~�M���z���a��F�m+�H���"3�������P���A��{=3�,�j�����PxY��:1
������"ؗ��9�;O2On~f	�d�j^4Ĺ�M�0��tƒb`�9_�f̕�Oa]մ=xk	`����|X��*	'䖯U�v���q��R �"��q���R�D�@� �VX�,��$�M��J�C�[�oG��H闫.�X�s�� ���"�d(�ٙ�"[�v�p�V�	s�R�йr]%�P�z���$6`*��dm[�k�.���O'��|�R0���$_�@ܴ����˖��CRP�t�UO�?��� ��Z\�,?L��� ��ʋ�Ѣ��n����ݡ��n{%��>G����P��(��@/j��\켳���&�@w��;�����X��P%>;�B�.�K�If�<V�6ʲ(�R��0�6��V=��w���&��{���.:*W�'�K�,f�^T7�����Ԩ[��V���̐[l�=��u�m��8�r!��O��g���NC��{�6�"[�%���j@`�	��W`����D��9��]��J~�AiA]��4��
*o��1�
���D+v��щP�q�7bTX�𼩗SI���e~.Ht~�<ǅ�%��g��<����J8�ܧ�ɔ�$���`���\�A~�&M���A���q@f�	����^C&�I��i(��ꖫ/�yЏ�	$�h'=��I:7p��$t�ṩ��1���}zT�vy�gH`�ð���.(��k��X@�F/N� �YB�6����2;���){~w\�s,ع��ssmws��Bƌ[�3N����JN.�SNa �薂J��3��}PL2��K�-&N���\<rS��e�O��� �d�~�ג�^�J�%�Z_�M��m�n�Ӹ�L`b~+��@�z���(�;��Õ�]M�75,`v����,_c�ݾ�Bgp\��)6��?��j��D���}���$IK��2�,c�z/X(�w;~��5��������W���
�ն ��[-+�sz(�7@�� *���r�Ol�ﺟ �� u�v�A��	�:T�B� j{�t"�{!��4���ڔ�G��9`ͣ2��&��H|.�E�ͣ�
��y��и:�>Z����N�:u��3��k]�c�^�D�$I�w
uӿU:է�G%�Jޏ��p�����(ǔ^�D;�ز���Q��ֶ���<.��j'h9��}AD�o6�:$��Mg�B�m0��e��\����!ۤ[� H2hȇl�<��%��TU�����f�ŞP���[��W���v��|i�؄�AE�䮔�($�����j|��3!�Z���6�y_w/Uo^�<^m$3�Eڎ�Y��O�X��n��Mv��2��F��s0I1e��Mހ�!�6D��*���*04�aQ�.�N�����۱���{l���'�	��PN�%1UF�?!��=���-dkr]�U
�bmE�p�1��4��k�vX��E<��E�B���Qw����@"=$���"1�|�<Ҋ�ЛRY��(�[��o�7�g]����F�W�:��<���E�5p�:�"_�Q-��[��ϡO����63l�����L��^c��ӕ�'�DY�� P��Z_\��uE����������AD�f�a�+֩�D��;��x���,��.�{ Н���<��#r��9q�;�E��������)��V�����:�sL��n�J���3�|�ou(�9
�k$�U��l���R�b�`r�i����y���!E�
�QEP��y����6S�n®��M�/��C�[�k�� �S�.%{��X�4�5k!� �?Ɉ^�I���$��h:�7&��ڱ`�z�!g�+��Dg'�_M�q��&�'a-��Z?���&�;aT/t�>#t������x�8��T9@n�O�����[��E�3ʈ�$5F��HYp���,|�|&#G�e����w46�@�׌%odBɇ=
�J��G������ڐzm�S�T\?B�I�9�UP�:���
	�
�o��b���+�s��_�X���A����O�^�K̷�ƻC�;oz�p �Y��UКH{�׹DIշ ����]�eRR�zf��Aب�d���n�J��5�U�I$롦G�At��p�rG��6O~.�p� �3c�B�K�h�g�9�,((X]��y��=����0�
�7�K��[�|5U�� LTT	�<~����J׼�".ɫ�_�Rj���z�n��B�Ek5V�B͢4Ȏ҄��ɼp�,� Y�Y"Hn���k�q��5>�
���SǨ�������FC������n%��� �N�r�ܥ�p�N�u�إ0������6�Ҽzy7�\ΰ�Ͻ�Z���1�Q*���B���#��.��^�t~�ѫ"������dɬ����|��♚K���bmZ�?Izb���ٯ�^��V���Õ{�I9:tO�Z@M4~ Hm��F�!t��8�H+N��Kt�[bF���{�!������:D�Dq/ޤ)4#P`\;���c�iM�M�]:�#k�gF.9�n����
�V\)u�M;�^nTZȖ��DwI����
�iq���NR��ޘ�D��ǉ��"ք��̬0A,�=�P��<�'���<�;J3���Xsg��f�܎��pj��\!���������}�)3z�[c�2�����/۟}>�[6C�uc�ٻ&��H�T��G�5a��̷A�`���6�$jR�U�eFpV<��r_yBg����$�m�=����CL�p�2w.��4|�r�l�'��=������D�$Q�C�7��r�֓���#��14�`�
 �K���c?�e��kз���o��u�|z�-�_8��"��b()��e�X[�)oӴd�lqn�'���AJ���W�5k�t#�'�A<��,��s7�a"ꄾ���.�`��75�����̞��~ڸ;ŝh��{���޷UT��.e�V��5�+3%i��R�2�%����XKY?��U�R�膩0�K���U
���Ղ&��A��n��w��̠E�S!;(b�i���b�_��Y	XP_�HCxA�M6[�Iؑ'���V��.
,g�
F�ש��8�B k�6���3�\����$AG�Xs0�)X	���#��C�R�����]Bzg���|T
uP��|�4���6�g�A���h9R3`�Nqec�ēy�xL�:��vF�KUl_0�t��y�n��(�o��Gi�]�=C�YIO��U�B�%թϖØr1��J��.M�1�o��ݑsaz�O�B����if%̳�׾ӊ T1���ʹ���Mu?$ M+��((�nHM������f����@+���a�"��3H��F㼇�|.�����t@3J��u����Vp�靆�k8=�SZ��t)��X��&n�+�ln�J���_�ׁ���YF���V�������	*��a�s#�C����<"�J�hVD��VS⁸ٕq��P٫��=xl֑��lk]�_.��3�/�\�qכ�,��B�wTU���9џ�|�#.��Y}�yS�p~J��D�g���G��'�z�Z�ҡ���B+���҄�6SX	�gd������~?*�ӇhL�Σ�8`��*��	���PM�ʩ�QN^�s"��㒴����] �-�/���OH�s�G�Q��p���G���W�|G?�(�8�sS$�,Q��"2�33��+x��$u|��e�I���[=ަ�q".�p��rH:�!��{�9d��z]7��d����W�4d9��L�RCh�	%�Y)��=\h�#o�p�U�����
@P�+T�Ҁ��+��=�1��
8���׌�m��'���Q�G����^|NMﰤ1�u�7v�/.�#�p&�Vw���"K����j�m-�z��@k��@��[(�������Q�D��
+6��{�����.���U�s� �2E�L&Q�A�yF@Y���Fc��>G�i��]����m�a7��[������hq�g��i>4r�}/=�@nϬ��@�=ٗfF��l#?S(�>#]b/t����T�	�-U2�ྑ�6��8Q|�<�s2�*k��1��Zf<_�ot��Ce,u����!f�.��x�*9nq8\�����������0{�~���da���(�;�S>R�V�,�����B>�dt��LΔ����k#�qV�&Tr˵�B�/%dPH.�[�ߝg(��k��H*@'�%`�E��Mxm���ٺ3��"����;���"k�Pd�փ{ms��g���(`�0���y����~��N��,��v�0�Q�!=cn������8������?xc$���&qk��/�zsu/)��j���"��^1uC>N�M�庸<���$�+2��������B������鎃�d/|��Lֿйy&�#X��[骕�;�1"�;��\��9�Ue���W�VFoρ��{�0�v�~@
C�z��*{G�iE$�4�\����f?�؈fb�ŘR���>�{/㻕{��YS���F�Os "�O!�*'��6#\� kJx�x��J����7�tӾ��M�2�I�	��L�XE���vl9CX�9�,�<�� \�����Ֆ��-/���as䭒6�������L���V�j,R�d�]�t�%[ľX�ۨPϊL`Y��FY��V&��eW��Ik��U���-�r6&u`��2��ף�{���
���N��+�Х�����AY���?���.��*Ed�������C��"�.N���얅ae�4���b����W�Bd�<�Ӡ��%3��dp)C�U������DF����2�*Y@��4t,t������Z�*�������H1�՗���C$PKp�ݏ��'�#�W<I���
��CB�� an��7�#�^�Df�B�����*�4`� �F���
;���yh�U�2w��I ��=�Zh=)s���?ծvP���0��J^�9��g���k����U�.�5�V���8�/�����h�-��I�,���/e�yC���0P��K?$�7�$>��R72�t8�G���/�&v"�.�ݕ�jϽ�|�t�O���}NW���ݙ�`�˭�tU�6Ǵgk����2��W$B�vwxwA�����/v|&li%D���Ĉ�7��Y�o�S����H������l�uW�\�k�	d���A>��L�5�|�j��K����/B�ofd�,X�`�fXu�-e���)�78M.��ESB����-�˄蔶� ����5K"��(op1h{�8�z��kK��<���A���a̋ŕ�ճp�N�c�:[B�>�`�5}���/�R{��q��+�F3s
����44��t�/�9�r�(����⩅G��R�ŖgI��JŇ�Kb
~i�w8���C"TlF/����)��/����H8^���,���ByM���lZ�&�Dk��/���c`�P��F�H'M�@>���Im#�K�T�(F�V���@�;>�?po���[x��<����D�*��a����l������	�UNr�~�f�INt�s����r�މ�b013��I��6r�ኛ̢�K�}	�o��U ��ϗ�1��2����P�$̃L� X8�Uvo�YF�"+��~�,� j��U���Q��$ԧDH�E0�ALI�3��������o�)=l�����h!.�&nv+�%��y]�[疬!� f�KHij��0�9Z�ߋƫ��q��Z��VJ���3.� �i���X����H�Ƴ�3A߮���Y��ų�}q%�_�{D~]$lN�a�F�yS�i�����2�=;��C�R��N>��DȲ�>�a={b�	b��"6/�OZ���.@�TdtN�~�B���� g28v�:|��-�a�xv@tV�ҙI�?�T0����\Se�����ΟP!l,H����J���bL8+q���0�10&f�s��uN^��}���nxƟ��[��R�l����0q��G_��� ot ������;�tׁZ2F��� v�!h��?��X��P������g��,SL��W)� �D׭�7V;Zwp�a���>�b�>o~��a*]iܵA�!9����������d�v�
��gnBo��8��g|S���ȑWA�d;��v����Ql�'�_O�����ޙQg�"�4^��}�㥶e�ȓw���PN��NFo�A�ʎ�M���L�����;�%�5��˸#{ؽ�FG��Ba���_��:��J�R�52s(Nf��.(�Ҕt����h��g�o�+�K�%dk�(�+B@��7�F�<_c���.���B%��@����捷�ȉ�^(��Z9̮���/�;�/z����vڡG������Jyd#�=�".��&�A��5(	6r�/{"ӣ�r+��@��7�0>2_}�FK�]]�\*�j;�����R�y=F��j�+'����:�Dd�8���1޿�Ѐџ�8a-�k|�MS�h���i�8 )p)�� �Ӆy��]ÿC�~WO�֋J��В���N��Rf��r���J�cJ �0+b	|a��сP��7*d:�@�h��o<���(�����&���N7lq(����l���{�H	^�
0)��u��ٻ�-A������-_7F!U5!�w'A�b�0�����Jc��5~r���.�&K�=�5g��΋�ؤ��0>>\��[&�xw/%���z��ve��9�lj�_���Q�',ؔ^-�O@
��v���� ���]} ��U��;!1p�&+�G�v�9U+X������V���H��C�0�F����:y��!�A��M�O#��וN����@�vv63��߸ޭ�mh^06��asj:�#���0�������f�h��("*$ZI=�}��qctc3<h�8w'���u�~�/��盚�9*G�����z�|�y�r�7�+�P������#0�;��~�4�k��Bbe�%�=�/_�J�8�;@"Y�i`���
�R�4�ʘ��7APfa�Tjr��پ!bq�m���y����KV���h�Y��kU]%�	�̹�
k�Mo�$����ƻjmE^/r*�W��������§��ɀ�NH�e��r.J�g��IN��1}�)��~��2��O`J���oUi���WT~�&�W1�+�����	�2��D�K=�
.T�ұ���{�%�4�G	�*d�o	?V��-�U�g:@��~}EF�c���:�Ŏ�'民5��� �m�P�k�/{�68�s2A���mj6y�
B.��m�J�%�:�l�=�ڹB{�S26�דvv�9D�i�Gh%�� E.,��C<*?����u�x�G�u��^��Q�:�Η?L�l�r-�Z��7z8ze~��\ݪ}�� �3��tA���2~��Vʭ�|�:��sCq�p=�@RC��u�����~�I�_�!|���
m��Uo�UP ���$��?c��M���!�d:'�1�u�����yjgv���"�۟O�\��� �rv�NДޒ�a@��[)!��ꔃ�o5�9�a%A�]%0�_��N�p�ϗ� T$Zi+��r�V,E@�ƛ�ˇ���6�M��hSO�Q%h�ܕxF�=m�G�=��1�E�Ľ�.���_sMx��${P3�U�t���V�Z\�1����G����* r,�/�6�Z�-��k/�ЩV�-˘+ C�	7U���Q�G�)��n��@�w��z�lZ�ʠ����H6�6�.��`�_�/ώTmqRQd�.F�-�N���t�}1�����7̯,��H�� ��2��rFo�'d��M��!n��pDvK�ҧ0,j[��P�~m�>W�x��δ_�aI�>L<q*�*�^��ߢ��u1��'2f��+��%lC��P>y�Wm�ѯ�6R���ٕ	:�l6Oo��U����5���ЍKV�rF��X)/`b��D=�1�~��ɝF~�SU%n�,w�-^v��8p�0�9��@!εN/�ΐG�Oe�A�g%�<q��I8q[�T���ֵ��C�cn(���,ɚ!�W��3��}E�~Ų$��F���*�|�5$�J�c�r���o�n
��\E�w�G��wӂ1(ݭg�P�;��o�,�yE�č^I7�.�.>���`ڽ�������\R�1����2���M��	X��9ș��x�T]��˴�Ϝ�m�l��_]�%ˏOݶ��d�BO��fd�q�-��!m �{`.������]L�m}��nub��/�whh�{K@iP��gފO��{���."YK߲�QQ�932�;c�}ڄ��q1htT.��"p0,�}��U�u{s��/�/x��s��&����_������G�O_�u4������(��b��%ڞA��ܤ�0��w�:��hAgL��Y5gu���|�zT�|�@\�XE8���/Dw�M� ���
͏1ֹ�鍱���-���?
������A�#	�����xͭ�����|�e����S�$���j��Z���46��1+x��3!��]�/�֏n�I�v?���P��I4[s鴷��}QK(��9ul�y�f+��!�<���eSJG�OJdL��9ܭ�\��2���.����9�8�|�#�ՓgW�ڮD��BFܿNt9�^P%�#g�z>�~�n�ѣ `�"�%��,?�E�]��:��O"����v�]�<�A�C<t�ݐD���%�fUT4�D�y�m,-q-Z�M&=5�=Z�s|n��6�p�0�^�D�G�ꗟ�$�-n:�<���w�4� �D�S��&r �ɉgK<_�[#ھ������]yr�������|����A��n��l��uIP���`A�V��u!���v�(�䇜XQG(3vt���Ġb��7�d����}+�	`���1i������Ӑ��������)�*?SbDX�V���˪���9ps�nE����2�uK�f�P�����{l���Te���������-isSu��\2��e��ɢ_���s�pGR���wK��ZxHb���BS������y��
��,�κ�"z�]즇Z����� ~X���z�����	�&�G�k��N�+��sYAn��#!̦�rk���uj�§༲x�t䥡D�8|yv,�`�R4/���D͸o�f��1��̘0��u2Oml�ܳ�O�O/�9q�����g���p�w�%�n+���6������}*��)�t�T�Ǫjq����KR��M#7��.fkAh�z�yj̍�O��b��=��3W|�
��l�̞ ��c~�0��������.	nX�{&#v��W1/r��藌�o�`Հ�Se��xV	���H���* �Bݿ�޴���>�=���\����ȅ�*��fq|�˴�Q���s�E
�ǯ$�X��l$7��E���1�K�mv���4�w�;Ĉ`�USW���/�?�4 �Ys�К��<崜8���^��`Z��+:��W]��ku͓���)�H���\�V'}���#���ӝ���#2�X�W��0�~��-�~i2k���_Eݪ����8��r�r�@_�1��NM�׭��QL�EPc-�XƅQ�j�4є���Ot�n;cr,%��>�ʡZu1k*�N�\�f쵩��� 7���WR)Σr��+�D3�-��� �X�#y���\=w�"w�(�8MLĘ�޺ �a��8��(	���3��i[�}GuJ7�����t��k�ɜ:�։��ě�Ú���PIߴIF��$+�I�}��}�#xE4z>�ĭBx�Av�S��V��ck�?��|3iB�+4��L��
Mx��a�U��i9�Αh!�)��Q�b0e{���YxB%SI �r2>"���Z���Ԝ���i�9���˃�#ŻXJ��&�Ù�"��牜����ت��D�����t���A���N�Co>�|�ߝL{U8P�nR���,1t��uٍx�ȸ��Rꏰ&84���_%n�0�F*6u=s�h�-?�x˚;�$�Qo��{�_���xSɄ�����t���K�㚝.Зb��+�	[��]L(��9f&-� B���-�ߌx�%����s@M����p�^�@���ޘ��l�	\�)9FJ;����X��	�7\�ݺs�6��[�轈��n�pk9�7ӄ�r�vՅ%�� �=	�5�}��IW���G�"'ҡ��+�����	ee8����3?���>��vc�L�����Z��'��'g�D��̱�0!{�cjW�K�0��ޮ���SR;���B���b��烈E�R�H�G��� $l7�1a�LL��_�HL��q�pa�٣$��������y��*��KվV�s6j�<�'�w�=^*ϥ� ��2i '���K��n��T�]U�qv���g�°Fr��?aXӔE�d��H�#`2�,��:�m�'h��Wz�{*M��6��+W�Z����;\�:�k��}N����nQ���_ֆ��Kh ����&o*%"^3B� �;�S﨡W�o��^�ш���Xj��N�t���^7�0��_|��*�QL�0;s�d�\?���C�z�c�t��N�J�qx>��K�V���r�����ٻL�9���X�ER�FG��w�Ҿ����̕!��.�8r:��^��͑N��޵%N3���G�<�76�3�e�������E�s**�;����"��������x�ˊì��(wc��Yv>I������~:}W�t�ޑ]��8��I���"!�W�O�/�V*��:@�����{S��Lq[h��������r��="b��NS!��i>
BYe��jaK�J%��%�tZ�OlrA`,w��5e��6�gԖ��n��@�4�ҋ�8�P�\C�h��;Lp~��Nu[N��C$���B�+`�2to�'����u軕~qK��Ѯ�������I�d�UwS��=X;5�y���X��1����qh|z4�Q���	ՉZ(��{��棅�K�Q���	4�Aʨə̥a)�]�1[�@��xț�x�*�'��v0y�o��C&7_q0�:޳�5�02���+aU���[�l}�R!��KL�݇Ӊ;ʪ�͎�TϮQ��xȓ2�0Gb����Fs=���P�Y
7:�g�\d�k��g��䏚����ySUF����t��"�%,:y�iT0�_ʙ�xGU)@�<r:�7-�'��L��m�S�z�O&z�'��KM,�9�`�{��p�b�[hu�h�G/��y�"D�Y���f��9(�Z`3��ȥt5d=G�%G1�5�<�aW�B���:����Ǣ
^�@ʑi%z�D�8`��X�C�����,$�� ��ͮ�!wx�����m�l'[���n����r��.D����4�1�-��?V�=1����l����6�5�����MO��E�`���-D�_s��YAI@�+t���$�h�#b����"8�}t��f %���MG�Q/(�7�8�٫��"���gmc��q%P�݈դ��#��h�e�.�@�S�h�GA �f:����#l�� v���Ե �p[��m��9�q��tyq��I��{����X�@�'�j?W(��ÀSY�u�B��m�E
�Ճ�[��mÕ-,���H��5��Y����6����J���B�7U��)�zh�	����Hv��̍+��=���s�R[���]GG�t� �ϴgA�[��YS�У�#��'��特��C������+^���i�?9o�!�l~����ݸrT�s�K6�l��T>����VK��]g�T�6�o-�1x��Jݣ�/�HZ�s�����FZ��x�.�^�$V* ��n��;�B/���mI��~�wP8��k⚛�U^�e����l��QO^�+�Dt���
��v�)~�����2�I��G�����i����&8���.�4�par���R;�S�m1�!�b
�	k�}}9�`����쁖�.�ߘ	�Ek��<��f=@�+C�RN�)����*ǀ����F&X�����GVVd=��a-Hٺ��_M(��Nó{�?1��HQCw�ٯ;��P��D�0�
-�"�)H�C������Рf�q���5������yփ�,-oloT�ոR}�ՠ5N�L+��񗿗�����i���#�`�l�[�x2F���k�$Ff}���5����!�;Bլ����HGX���C��/�,��7G�!��#��n���ZS�w%i��EQ�_��r�\.�b�{\w�v��_'vLғw���a�e/�ƍ�������ɒ]���5�hv{	*,x�V$a��H�E
'��E*���b7Ʈ4��Z{�NA	�I��q;t��;i��m-�̾�I�(���ØQ���`�����[E��17a�

J�#)ܷr�s���o�|J߬���~����\x&�n��gX|�����;�,v"FD�~�G��g6#9
s9������aތ��Ե��H���b���p���0�|2�;J��'b?�`�_�6SЂm�D�
�S�y�ǐ�����@���R���}���'��<$�֥��5�^-9ޭ��/K��&5I.�D��}x�{�0v��^�?�_�_�I����G��K~�O���!��	K�Do�
M�_lLr*�;gh�
@����єtQ2Dc�J$P���)�bc�K��N�EF��6�D����N���Vת��<]oY@����q(�u|�ߎg����-Kz�[�L����	��A����p�4�夡�$Uިu�h�ET�����^[l�hؑp�t���X�w�d[߳��&:��Q��)/���0NkQ�sø��+��Q!1�^&ƠZ2�6�7PD�?�i��>�JV��V0ˢ�S����~�S���U�%��2qS���k�I�������l�QG&���C�ƕ��,�ʻGr'���E����'f���l����U��t �]��Ig�!�'*݅a��� �
�H�� ƹ����r�0_	E��6+[���&�2Ƒ�r���!%]��kc�FQ���*���N�b'b��]Hu�	��?���s������˹���m�h,>��s��nFfS�q���k���~�9l��L}I�hd[?H���e���QZ�� >����Fsa�ur "����̓��I󘪴�D�|6��$�	�Z��z����w����ﶦ_�Y�$����~�@(��z�o��@��F���(�+���т�h�đ��ܒS���Z�bCWfd����:��4��$�hD����c�ۣ��*��]�o�q3j�B�Z�b�� ��xl0B0"NvY�/h��3&�FPe��|�>�kԝ�+�M��\�̤�U)n��Հ3���3ì����4y���F�g©}�NO�RA�CG���l޷ir9�N�Z�HO;� d�>A�32����Q����-Y[��U*S}����P��M 9T&�bq�C�i��WBܱ� ɯD��[�Dq�g���/�J��ĕ�
M���f��νĒ�)٪}Rj�b��V���E�fiN|�m_�����Ễs}y]ѻ$��K�w�|w%[0	 �]ww��'ْ�&����7[��P}z6��Q׳ ò�MC-*Bsr�L��q����E��v ���d�E�h�0��z�ӉT�
�0�T[�l8�h%ĝ���
�U ׈�[ǅ���b�Ct�v0�D�Y���.�S9G;hF=/��&^ȍu�lg�� 9��5���5���c�ճ�8�V5��i?)w5��l�ǭ�K��#���ZZB+�.�ˍ�9�]���8
>��ɑ�|<����� � Ʒ���̔5�X� #ki5�/�&����>�\���Q?���p�ꥒEX ́e�C�5��eu���z��c��5I47MѲ���["�&�p7�>P�7o,s�}�JN��bS�,�g�uԔ߮�G��o��a��m{c�'p��_W�;X>�X؁-���U�P�w��u��k&���@���P�� ́�Zb�7'i��oW��Ƞ� �6�OD���_D�=�np�^�TT	p_IŖ���9P빨�7��M�J�r�ǟ+V��{'4��(e�a���~�
v��\ʖy�/�v�~pO�H�>��P6H!^�IK-<�H�ad������R�u��-�
�dW���Bdޝ��C�E�l=ܤ���?��P�巷�a���YQ:j�\�,�F�EA���re��81=�/O֏��x/��&�>S9��|wI
8Ha�~��Ċ']���c�F-�����+S�'�����Gc�A��j��b����+e�U!�<�&��r�ԍ��?�*�mLn]���fWq+B�2�	Co�8 �D��$E��	L�&7����%����)�};V�#�`k�{[�T��D˻�T�]}��5�����lZ䧃v:�A�������pG���(��H���Cf��ݮ�-�4���E����ky6R��ϪBkx3��F�՚�ac���k�R�S�(�k����Iˤ�d�A*wA]	��#�}L4�� z�	��k��hђ�r���g�^0��D��;e��X���m��;�<�l�:��ܪ��XV���E8�de#�Ƭ�{-����K�7����Q��b���A�L�IU�a��\�ɶ~'"q�9I��琛aڡ��zx�	�Vb�gx�9����7�v_���w	���2��_���l!]�|�;��@ gxsU�X�y5Ċ��#6�-�����d<|�i�������P.�KP?�tJ-��PY�X�9���.�YT�r�$�c��Щ�j����Fd��fN�_���?�Y��ｌ��ERm.���2_Ӏ��/���ៗ�`����ճ��5���.�NP湏��,a��U!�,�9�Eo���s� �,��1Yo���D�<(.3�#�� �䨼: 5wpUN���A-���ڜ���]��ל��H��ls����;l�	��;2���y���i� ��v�ص��]GK���x��{���u�rC2ۓ/XD����M�u6�a7�)�cyn����c�Y��&��ͦ#�y�ygO�~qO4$���(��U�v��f�����,�5�ab��;���u��$��Xr��h4�/�@X9@���?>�/��~��&��JU0۾l���,��p
���s��|�p����Rl�;8�4����աy�A�[C� ����ǖ�lz�q��6������#D�LG)�����^�qX��"�cG� 6�\&�g�D����P캣��Ik갰�0,6���Ė�vJ���v��ݏ�`dt��o?|���:���e��B�F~�'Jiׂ����]��?>�z���A�5�!�X��Y�Y�A���]��ʘ�v�+�ob��Ϗ���K6���Za��ļ��zo���P�uP�lP�drg)�]�o��d�%Gn�q�z>�&ٵ[I�V�F���K>������ �v�GǺ�K�^K`��'w?��Z�/r̍~�G��$�qC��2����c��1�f�]�*��6p�@7�E�<�d�f����q�xqMD��O��4���MM{����Gv�
J��5~i�P.�p��)�N�'3�b6 ���}�)˸_tO�(��7�h <����ьɞw0Y��Kv?�b�A��]�%>_g�n�X"Ge��9����r���Y�@�L���7d��iV-L�k�X�G:���1�%j���}����	�7��B,��^��}6��]8��O��Q�qL�1�J���=�3ɣ+7)�/�����H��ĕ�|BB�ߓcyX�+�)P�Ⱦ�����1���kj~,�\/��LP�H����-b�8m��9b[������?��B(��6r�P�o�#��4��g�'�����Se+���	�~tA>"��9psT���GY���΀���f6 ����cH@�?Hp���v\*�~��]G��8�Q;�r<ng~�Yx�-�ߦF�|[ٵ)x�XS�<�i�~�y�lZ�d�o�X��$�3P!E��r�̫�1��@�����[p�P��wB��Q̋�S�����&�0Nh�Y�?`�6)�x��,cB��XeKf��y�}@��0����o  �C��$�$ʡ��|'>49�]{Wʶ�a/F�*�$���D`4��q�J�\Z愩��3�����#�	� �H(��̒�$�� �a��D_2�@���.�h�N�ᣏ��	g���\��]q?2�1g��Ǒ�(�p�g��r�r�}2��rg��ѿ�P�y㞫�;LJt M�<͌�� �E���=ޕ��:4\�P�"W؞߹R)���8
�4�R����
-�E��+�Ϗ���9ʦ�A�T�qa�lʍ�9O�c��y.�_��&3�D�bw�!K1D�NS]urp�,BpI⬠�AKV��!�O�4�M�p��T��r/x�m2�7]�.^�Ec)+��{ y�j��m��TZ�L/G�Й��d�Y�N(�Ќ7�8�^�%�Ԇ�[�xG$톗������B7�cu_�sx��k.�{�ê�Cm1�Ó�g��ݶ��@S�� e�+���� aY��n
4���n=4C��AY����f��<���3�C�M`�_!�������)l�W�*��f<k��CDW�O�i�i�2#��)ǖ ��l>�;5.�������Wɹ3��H���Ԩ��`�g�t���;a�y�+�2*�n�ذ��F�}Z`H��h�"w�$���0�.Q�I�=��>2O~�3%�bo��אJ+'���ؖX���ͩ��������䳘�@�Q� 
H�����ㅪz#��+>$*�nyk�H�?j�O�	L$w�u���M���Y���		�y� �MoŒ�H�A --nL�zbY�~�R�(�\��ZG]��C�]�0EŨ�!~�R�fQ��M���R�s4���7εxD�x���ͭ�����c<�����cjM�����X���I�i/TW����/x9���d��y�N�۾y�
I�+�	<L]^��6e�{�x�y���N*4*sM�BR'm�|I�j��ן���:7�_�K��Q�v�r��-J�9ݺ�\w6�[n3r_A^{��*wp�[�Эyz��^�dէe!����:=l�s8���(/�u���$��4Y�k
�@)�_�<Á
+�^�2�-�wQ��Խ�&���Ϋ	�"��H�1�i�kvz��*�5����U�	�1嬘�S$�um�TF���8�:�a�G�øm���?��w`ʚR�0E�X�����7GӚc	��q�p:��,��W�g�0��F�p#c	���p>O@{ڀP>�!j�^'���3y�oS8��ꨴ���%�8��e3�c�� Yw�Q� +a�>Cu�)�r@�J�_dj�Ǹ���=o���;��oD��4����dZ�l�a?eąe����9
�;�}ӳ�I�ΤȀk�BfEh���cAcn ez8�J�+�倁�t5�U�P��%�+V�!�UV͍�o��v���݉u�#���ȼ�� Բ|I]��|5�''ݲ���-w�aޟ[CC�1�Wy�\J�J�.o��P�	$�yA])���'�f�F	
�^I�)��M,���d�][����0"���m,i����Ԧm4�]��YfO;#)�{��7��6.�'Zs�K���moi�_Dnu�gy�६r�u����$g9b>hf�SZ��S=�$�c�D`������7���R&�j�`�|2��R��~@Wd�u�>�GP'����S�DO�AvĆ9�\��:\��@�އ�ɲ���7\Wx4'��V@㥖�g%�u�#�o��{�ulߕ�f��X.��O���X�!\�@Ά.5�a�5�L���
��Ω�hr��N����N��=���_T�y�ČZ�BO�b���p�k�-�[g	���C'�KHP* 覄dڶ�O�x$h��A?����M�-��gI2��Sף������UOc��F搴LR�5��xt9o��zOh�ު���
�¡��?#�jufo�hx��cA��,�j�Al���<\&�<)&^HR�����b��y{��8�^Ï��Ƥ.��|71�C�9��?	���n"�a�/B�W���M���o�v)��5�e�x�8f��u�p�w�"n�~�"V�_�)�ы�с}	�D�x��9��<@�n6��ǞHv�m_��������}�s�F��]�k���(�T��E�*<ؒ�?���/'QM���X�F6fwH�B�%n� ��3$�K�:I������}v���|�hN'ZB��*;R�?	��4��s��X�sG о�����IOEKغ�eTP���+�}��Еޯ��o�/9�H6N�CO>�W�ܘ��H�C��B˲a+�����^�9��ʈ��l���dP��|.�� [Ђ���Ew>�PY�e�����`fO�n����_������&� �~���vXA�|.ńJ����͔ր�1:���3�_�US<�Q�w[�:un:|wL��g��Z�_;��T��O�}��A�*�\l�����$�;\��TCs"�y��>+���@XS��L]��B`n0�u�p�?�gx�b��  g����;�H��_m8ܬ�~Glb$#;�#L)�5-9'AV��/K�#�b�b1�yľV��\�5��5��2�v�W:ц��C���L�72�TK#�ʎ8Λ����%��* �@��(M � ����cI������w�w�|���^��[t��0�9�~W��_������\�@	�L�������Q��w���u���hw�ãI���5�k�L`1�ժF:�Xg�l� L�7�*Un{[�, '&"ɽ�l�3iP, �����`�C��[��)��6��e�]S�$�fJp�D��Q�Tvm�y�t^G������� �q�d�`�� ����

@xM�g(�D~84WC2bA������1���.	�&�F�z%�3[x����*�y���v\��}���_�蟗@��n�Gd�.],�x$�u"��6�UGs��
s�S,����y�����a�O/�a�<�By��m�k>ѱ�,�
�`!d:��tU�J���N�Sh�J[~�����>��_�Dػ�N�9�����u�����w���wh	��T7�r�k��n/\��}����[o�"�g�����<�� �$�Sm��3��B�p��v��ه��a
�[���,z!n���ރsY����i %;0 �f95��l%j��6�]��췰�XzXJ���_�����TU���7L�#F�����lѹ�r,�@J�\p����L'u�<������%x�����*�a�~�����o�����@�z2%y9q\V[���GHUgUc���Ώ]bLЯݰ\�1�m��_%�&�.x>u������v�Ӆ�H��^t���o,���ٝ��Wʨ|�+T)���J�^��U�5��
"'K}S��*ţ2���C�`1ί6��ZBv���G;�p��wx�x_���0�lR����K7�$�T�Ul�-��ߺު�v1�����a���6�������{M����ɬ�c�?��^񼟝<G��BLD4�
8b����k�c�PA?��K���?��b�1?�"d9�F�g���ۃ.�� �I8훖hc�,�#=bl���2i虜G�$=S�y¾�.�tç��_���i���wмJ��1ՠ$�􋭁z�Md�~�;��j@��5`�Ɍ�y7_0�y#*�*�j|��	7Jsw�S�@��&VMӅ� �d�/Z���S���2	�������K`��ra��Ȋ�G�����T��C決�:���%L�GC£��"3��M�z��)za	&@E=�X��	!��1_�NZlq"�W�h�ݶU��MK��{)�g�8�w���ϫL��%�QTu�q�Lַ�b�j*N:��_ҷL��"���qޯ49�_�w���m��_�>���XǾ�7��3�%���)/.P�u��>MuD��<pq[�d���2�6��+�??�O�^*�����tF87Լa�>[�?|�@�K��7�pm�`m�%/my{��$	��QBfc�1+_�Gɡ�Kt ��"�0\���?%Q���VoO���d&pK�P�x&(�Ŧ�@�a믙д����-Tڙ8f���7�����9$����7��m�`v�����{�/(����A��=���}�c�[�?���c�B9sJ��e�U�F�.@�%�cD9���zqe �h�ʶ2o�m�"��|�����%�}/��U���/zs��� ����5!����h�C��������eI��7�I>�a������������*f�H��rV'��Dí5�	��'���R%�8-��k��d5��w�4��t��,�_�MK�V��0B���G��RZ�)zOWy�j>a��]� �L�.��Sfx��?ӣwV9�u��.m�7l7�Ɩ�WƲJm��dL����{��,/�����m8���Y�&K��4=�Z���Y$a
E���}�D3&M����Ƙ�Ϟ�5��A/�lV$#S�#݌�\~!M��I;�>��$_���K�����;�g!��C���7������*.;N��I�\�⁆=��%� �"]���Z�LP'5��i��CQ�+�4���]�z$ƵmV��#n~���.sy�� P��SY��LQ�Q�+�X+r�|�� �9
���3c���|sYh`��A�J���b$���q�F���%���4�ҧv��ظ��u/��+��s/,Y�� ��w�< Ů^S������X�|�7e�Jtl?#p��(PJOO��#��q^*H�����WS,��D�D ��R�~���F6A���2E��јg�4O�V|"��8.�d����B�z�Y�~�\j�L^t8�Q��&�������y�����<��iD�U&Y��e�{�����!�r��5b�)��@�x=���@Ҝ��;Ac��_�c��?<u!��P�f�E[�#Y�1��@�Oܿq�96 ���a\��c�l�o�(�=�v���)�C*���blw���k�EB��/�y(��&�C9��J�}�Տ�v����@��ȼ�ñ�C���s��*������a�6w�_e�YPQ��
�f���L\��U�8y8|����BԮ�.8g�B�IC�4l.K�;�u����+�����1�?-��T��r�{(�LO���`�Б���QT(1�ٶ��ך�h2[�k�}�)�%w8W�6L⾐m:�@ �$�y���8���J�5�
��+���S�z=n>��?�"�S{ݜ����5����#��HLZ -l���o�_2ك�';�%_@��F�f)��Y����f� �R[~?��eNH����A�7��L������*]d���ݐ�5&���U���B�$�@��r�-�+�i�\�ET6�Ϫ�v���B]��o���\]#:iN�����8Z��{��x@s�3]�w2��.�W|aCؘqPr�"��W���{���[̽`~�����IX��(���#�"=���Ml�ZQ?��v�O$��G�YG�A..p���'���c��xC'�+���_�~͇W�ڣM.rmf��m:�TOJ���cջ+[�)l�B	-b2�C1�"T_� �ND�a�㒿�X�ӏ`���mZ�Xt�֒4��~���x� �R�MK1
~u�@�0���X������i��|��+�1������v�3%�������Ƅ�ҸK�?������W�:��%u��3������T�Z�c�s{��7#yL�ܴ��������d��A�.&���E�t�����<�r�~0"���g�H'n ̬�g#`�`�"u��)�c���RO!���kh.��)+�_=`�k���P����n��XO���Y܎���]���Fh6��O�
���:��a�n���W9dW;Qv�}�M��O,"�^� �׎���t���KUdCU��'��o�n�y%lE	�`$zj)�钔)MD��?=�������y٧gm������