��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����� ����m��Q�D{S���;��ie�9ߧ)������o�A������5�XY�_{H�'�'�	m}u�QV���W�C�H�M���儙�.?T\���ۢm�������|湌�#���Y/.�W$e{�Y�	���O��K��l�b l��~�9��b�� %惦v��TtJ֝q�'-���cX���`�d��ƫ{���~�D\��0��P����o����O����B`)R���)��]XFjh�ݸ���"��������� bZ��3]�C>2�-p����Ԯy#ʖxU��4���!��U�]Lz�7<�`E���X�|�����;��:��/|����U4:�W�2�u��B�z$n�x�7-*T������S�"�N"T������2^:ofJJ�%��0��}�s��'�sرR"q�3��~�I�%�Y��R��m�"])e����q��=�s�w�w�TG�E?%J�!ju�@�NuJ�;��&�$Wo�^_��N���:���6��yU�i�vS���L�p�?+��F|��Ա�)U�����|"戍���r�vZ���f��E�O~\���|Xn19�C@�x%���La��
��*�(
���o���$_jȥ>J\t�^���[W��0A�|�0����*m%��L� ��}�1��@�ę�7�}����4�@d߲�	�w(���=c=$(B#��'̍�Q�S�9�-�x�N�W!�]��I9��5PmQ$�:�V��Gq��������xR*��|��)9�2T�krJ ���0�1�׺��O�D��8e�L��?4�)(�]��7�*k��;��Z+����&L���˞�Y�c!�����:<8�a�?�'�0xh���Y�0����'-��#�%�esn=3RYcQL&!�M
>�D5Lt���K-S{񭵽BN4���3`��w:��^��K�+�t�T��w9(����('ٚ����{n��haG:�up�W��R�4�j~�HN�eUiwą|�T�g�����dx�E{��sbb��o��h_A��lb����'�H�Q�u���.J��xC=��3U�;����}�����9�f�aO�5"�1�*h-�i�lg�9ub��4hҒ�T��w|[�%��/�� ��Ǯ��HɒS;�$C`H��!������8H���_E�;Ԕ_�4����3]9OMk`٢<�䘪~�j��3�d���U/-�Οi���s�_��)��Y4Y�k(�3��{]�^U<K�7%g]������#�N9�3{����������cҮI�z��uDqR4��Z ����J�[u9�E	�ˬa z��fƦ{1IU�>i�M+3 �`�`.T��q�6	����6c��}���h�*��㉙��x��q;J>�.@T��Nϣς_�$m��:/�'�.C�%�����,��ZC��: �ܦw���H�X�3�7���a�)Ê��v)i�)s���G�������R	U
�!88�[�A30aj8���Ζ܆Ln�o��Q����]��T�`�Ta�U�Gք�9fG���w�	�1�pm�I�*-	�)��e��isN��1~��m�
R��z�F�^�5�0odb>�O�o)&B��Y�U��¹���LI'��&ֹ��h��z寮Z޶DQJ��%�s��1�3����)?��[�����1H�!�KE�/}c��9�y��i��G=��YƎ��D%���U%)�.��N�j���ȞW\��%�"!|x��ʍ��M8���G��[���¥��h���zE]b��"�ol������q{���UO��f{�)��]�Qk�������o��<��n���\n!���yQ6eL��臤1oL�`LA�LC�����)�,/z%��u4�
������>�ŷHc�I(��Ws�?$�Z(e��"�<F{H5`�)��:}�W����dp��e���	hT@,�� �b~���%.�U���q�9�C޽��u�5۸���QM�A�*s/W�2An��/�ѱ�
oe`��O�!q���9;�y'��w��XxW>["Fղ�Z\o��|B�O�'��I��݂�b�
	 ?�I$)���֧���`��­|��̾�ҫ/�E�y
6�@��]��z*(x/�i��{���YN�� Oɦ�)���X���]�W(�_f���/_�NuE�20���B6���LBh�^�� f����	��1B~}�9��;�:�kNk����d����2 
 ���#�rZf�4���c+�������M��Ŕ	#����ѴKx %�w�Ӕ�l���ؐ�_�W����� ).�m��U/W�9{m��q��iZ/ی��!����M�Iu��zC��\bFX���L6���4Z�����7����Gl��Uh�v�v�\�7{��!]&����m8�NUW��Y��
��c7�2&`�"E`U�Z�붽��H�F��A��?�8]��d��qb�	�y�6
U�=!�W�UQ�g,%��[��9��$$8e�Ϋe	�Dd�oEe-a�����ﰌ'u �����64��{.�
]�'�i惞@\�M���oڡM��	�F������� 4�OB����Ɗ?P%����R�'P+�Jǂ�g�+!���šDd��d'���!m0;5G�(�P^��;8wS��e�y�ժP�w�r!�������X�HLH�\�Wݓ�>J������O�7D���I�����bglн� ��;�>�J`�n?#��E0Wf�H���r���r_+���,DZ���B���,�#�+��3B	c�КY���#�1$)ݰ����P��z���g��8-���#�$l���;��:��nz��(`�)�א>{+��3ZUu۩����|c����,�+�������"���	uQ�ݵ���(�U�b����+�'�t����� �vJ9�ô����`}y�j�g��j6�l����7�N����R���� \�Q>�h�zi��낱��h���z�Qv�&�8�T�m��߱Kȑ����<�������FK�j���:6�_��#��IZG��.(��Z�9JZ�~
�84_,|i��J���N*T��0��i�hQ�?v�� "ԉ9n�7d���� Q��
@jlS�T܊� _�L�*������M���gT�*�j�s�l+oX/���x��JYa5]ܤ��2y�l+<��/���qwՖ��,��u]�9c}��ں��(���+첂QAn�r#�<��
'��Ѕ)oG'3�==��[t���"8<�Q�sɴ��<�=VG2\�+��m�wh�[���6��A�萎����*|�ai�&���̸�+�kmb�q|bN�3�կ�0>����k����[HC��i����Y�.�����3�(�눓�6����z�:��Z��:��O���;����$�D��S�
g�׃ �l/�<���O/N�N;��#���F��������ŕ�b"[P[~]�����8��v�xt$��ɝz	rW�B��&Ǧ(D����[������ǟ�🏉x�"�J��כ��y��](�� ��?�����ؼr�$��6�� :ܷ��{*���]�p�=_H��g(�a�}HXnB�K��F �Ȼ.�@�1��=����3�Qo��qR���ŔL��X�����6bk#N!c|���
�4��d��W���Z�ӒP�>�UG�'�f����c���B�$��:�z<l���pc���lt;jI�����Tr*��<�3�_����4����<�\GU�D�:"���x}�C�{_��Z_�_�w!�s���D!ֽwQ�Bk��s�6��&�u����!v��~��G:���0vTУ�- ]��݃��l_z�#�/'�#�K�|�E��Cb�VBW�x���c@���=�+�pJ��r*�e�[b%`/��!*ts�!e'ln�$���_��b����Ų�I<�ަ��?��Qj��7��PB����G���\�Wݎ�L=���9�e�K�Y̙��0S+�!�s�]�)�Ul�Q����$D�l���ȬC�
Ӆ��)X����J S@�򚮹-���'���/�cfW��6�'�6��樵�_݇w���.�Q6�M���<��ֽ�p���z���u��&5Z�ƿFҋ:g���(��x�e	�\����Ad�v3�!�[����M&�\�C8̥�4�i#�˘����Bٓ�B4�a@0ܵr8kQ6���]^�\7ن2����5��u�?i� *li9n�?�,��ƶ��@�}���UǊ���)��v�ڊQ:;��B�Y�N��:�Nj�\I�@^������/��S��ïnۦ�(~T���������T�����6�5/\O<J��;:fo��|Ԩ��E�%!� iw�t;�-��O�H��8���aI�P?#O]��=���ؠ��[#�rg���|��"0�%�8��@5X�@�Ă��f/S��G�i'ke�_"�����nQ�R8"�*� 94��� �F�0X63YJL�\Ğ��x��8)�-�cγ��tl��B�l����t����Ɣ�/b�0E�AJ�X�{d�e#o[�l��
d�3�!-!E%�+n�sg}O�t� p��~K~Z�FS�.�@ה2���ZtZ��6��3��'���p��gn�y)�H����7"Z4%��K���o�@ֵDL>!䯭�j�ƅ��.E��a.84��o�C�If�UK���j���6�o��޶3,_X* <��y��X����{�w��w�c�Q�M4I!�3����R#]��^�{��T0��TUM�ѹt�XV��w�+MwQk�
T��S�z��F !�y��0���ě3Lv��/��Ea�OR"�Q�բ0��^�H )�c2F�Do���E�SU:~�Tz�����z�b�W�z^�hT=!�z�����^�3*�508�<�Wl~,����E��I,�fO� ����X�<���
A�A���	��B� 2�C�R{y�{�,�&���Ы��+3�T���Q.VF֔�n˾�	�v�]�論f�������9�x�:��^��^⽇|Nȑ�:��޹�vJ1lr#6����7ݧ��&��j)�+C�8e�O�L[��}b�Z���~N�L�%Y~�F!�?D�f�n��R���h��9�I����v�V��/�/=E�C�+�D�Ր;b�� �M�kd��ݴʧ6�S����t��>�m4�-�T����5+���m$�ӆ��W��G�3_�PP-�W̢X��5�J!R�
�Ekh _����!��J/@!�ei��V����:��L��MTz�wI�@�[�������,�������v6�N+�LNr�.]��E{r=ɰ֦>2?eI�1��,U|Jٔ0�ȃ��{��c�	��4�ڞ�K����I7<S����3���}D��
�����y'L��A�DL���Dڄs��r�P��]~���������9��2k mX�r�m)�vq9L�������[x��<>2��L��n�9�����KK��=��;�ASt�a��o�O�!aR2mXC�X�K?�,xLh���S~&T��-&Gʅ�Sd��;���������I;)�����r6��׉�>U��^��@>[��+�Ї�鱣Ǿ�����U�J�/�h2Sn$ǳ�ret�cduB*2�9���@�8�ۚ�������mދ�,�^_���"��)
	}4Z'_g��������C���Ȳxn{��?{?�lA�����)��y>MP���ld�M��	,���pf�/�g��9!�bg���u+�?u�Ε�[b��jV	��u dΐj*�%.e=�!$+lD�z�x-ʹM�HbԎ[ƞL@�>�X`��9�a��bj�{e��AٶV�87s�Ծic����l���/�K���,��A���M�J��qc�WGifsw�IMۘō@�yp8�ml=�yy<R�G8�g���^O�h��)1�����������yo�/��i��Y>�6��g�+	�P����|���lj�j�{Ǘ���l^K~���Ζ}�ʀ�r
��Ƹ�i�`�����h1a[����q�m	���1�������\��좋�.'4c��3J<W��!6Q����S^$pUOb��������軅�h� <O�{@s�;�!ӎІf�/{ce�yM�������z�/M����qm;ÿȏ�`�5ZI�38]1b�B�CR8h$�����n�f��E�����5a&\Âx�����,:���K�ɵ���<����R����δ�"ۈ�	��sq���t�q�'�Ɉ�~T�]��d4�>m���zz@�����됇�I>��ӧM]�7���;��x��h���1^��C��KXA�kU��@3Q����z�Heb@M�s��1�Vb� *��J�����⋛��B��t-]��m��D��Eᖳ�0����kyN��}��ғ32F�}�+b��$�2�d{���/[uC���R)>b&JczԜ��
2x=Np�Uk"��Wu?�
��EY`�8��Y������sh<;߁��2�Y�S�iT&�5�"5|��S1��,�:��	D7��'#?`@�cv1vۛ�r#�������cg8{c"�5�Ñ8��-?��p���S@t��T�nsW^^e����%�c �ZSv��Ƹ�D�BqC��گR���U�x��of6����f<��82�&}�R��\����+x��QA�,6(�f����&�>ewuq�J�������;�;����:�;�����Ra�L�-���c���us0��X��<�%�2
�&��!���*��n&\�5�W0ē�&�z+����,�Py��s6��|An�;v4�A��Rѩ)��z2�=��ba�@`ғF�����w��[���g��V�y��k��*�����o����S����F�Mـ�Լ����{�?H��.�k� �`�����.g�*3���~��񼶐�Tq��{�eyÂ*r�-ޮr~~Xك[�\P�\p��2�h�z�XP�6 ��n��G�;7c]�j������1���p>���A�y,��pf��T��g+EITN糙�m��}�\.�o��*lF�)�Zѽ.��QE-%��
Nv	*~~8��H��+N<���fV�0Nt�:.��׽-ȋPl�����56Q/<:B��0c'@���W[6"���XO��GB^����MˢdZˌ)��>����_}�lF.(�O3%��ͬ�gj݄���=(D+v�u�=-�X��G�qmG��"�!�[���N�\��z-\���8tQOӇ�{v�d4M2N;�0H���P.}�%q)�R9U!!m�B`Y*y'A��)�lЉ`I�'Wo 
��	�'K��/4+�DZ8���`]��ѫ�5�k���>���g��6h�U[�^��Hz�8b����.���k��� � 9�]iM��@�a��a>/p�x8�Mۉجa�9�׏m|ԕ�a+3����\	48�G�q�%I�`�L[L6��2�`��b��gw��aה�����!9�Y��ڗm���8-@R��lg̭	ڂ<�_ p;