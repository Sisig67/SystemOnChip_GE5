��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%���J�(J�D5`��U4�(��c�/�k��iJ�(z�����A��A%n�YC��U�!K+�P���G�1E�Ƣ���S�H��ZkCQb��Mbu[ϔ�Hw�;��S� ^p R.���첗� ��������vN���s�\{z	�{&����4!u��~��?/R��Ț��9��,ds���eG��g�%R�VQ�w$�� Gж�>�33���*�ڭ�3���E��њ��b3�UL'��x�_P�A���ņ� g�h�ç�i���P��o�@O�xl�с�.�zz�f���F=����k�a*�����2��/=b����!�Ϗ^���%#Pn�ު�F6��J��٨�'M�Fn�^��4	�ᘾ�k��N:m�	M���s�u��u���dץa���}��d� 'W)=���eR��� J����F�03HgQ:}U;�"�>�=rMEM|�$�Q�lXA��N��$��<��A��Z% ={��)=���i��h���jl�ϰn�2��
9�O�:\�T��?\޿=�^_^��o�{�7��e�8�ab�x�S���m0���w~�
,FAI5gP�h\��F7��-�g|��e�X)� ����uH(i��׵�\d�#dH�,�+��e�͉mEG5_�z]�>���dL������=T!�6m�)gɥ�B`ܭA2��EbC�CA_�2��6���Uf~0L��;�#b�1�_.kA'?�w頨!�'ݝ���5�UWRt�w+"!�c�!~QQ�As8a�c˝*��@kYk=�5TҐ��W��Y�(��K� �Y�	����K1�2�G �"����O��Prq������#�Қ2���=k����Fت5N'i(���	�"�Pr9��X�
��>-z^QP�v�g�8(0b��=��։���S��\D�b�E̤���������F��q
bŏ�+ed�����;_�b��v��cH����o�?��eb-���8���-���Oj�O]ZT��ō� ��`�9�����֊�����
�G]CU�b6ȇ�f|��R� ���ޏ����cG�++����A3�I�4����g�!4�әB���5�P���/ñ��SS8�28R��Pxb�:x��w���I7	�}��<%���ͺ�Dƍp9�	�� _��Y���UE�"Qb��n��Ll5�	̼�b�/ �U���@�R~86���
I>��^nL�ɨ`+��4f�*#�p6�&�p�Ye`�t�,�
�V~fl	mK�=���`�5���Ls5���t�A�{el��z��I}([��{�|_���V9���#���nBt��8 _kk���z�X�ɧ+�m�B�����'��/l�5��W�r�?k�����c`ۺ�au7+�
�{���U�?1m���'�H�3)o7�&�b�v:��绑Jh���:�㛜�x$�y�4�Y�Cn�ף&.G+�C!W�$T��/Y|��e?f���!Q��x�������2^���<\��^��v�P����R/�|<uݲ�h�r�B:V���rA47�3~D�B��4�$��=�����h����R�x�f��Qh�亮,߀�<p!..q�N���Щ�~U������N�� G�l+iu�ÆXX�V�4��)(��j����v_5bM��Ϸ	*ڀ�F���:c\h�^d��ݚ`R ޟ�]O�%�.�<�8g��읟pQ"�u(}����2q~�yeL2`��h%7��9�^<>hY[s�[�c���u�;nS���M���"�2=���Mk1RS;1C��0̝����#�����ʂEU't,�j� au�M�4'0&Q"�<�����漶�����h������OQY
1��tS��R͆AQ�N�|E2����@" sZ�0mV�_�����r���
3oL���0�����r�<O�+[hed��i���r1�#`��p+#�5��6�@b���";��"|0�N�n��H�ν�bV���=�34���R��F>\����,ְ���ν�d�骫p����^����B��-�T�pX�v˻P�.����lr�&3����FRӚ)nb,����H��~3L~�Iz~�YC����?�I ��)�3�? siX
���[6X�Z�|�/|.�k��aG&,�|k%�Zzkh؃U=��^MV�����d��5F�&9u�8�Q��ٹI�AZ����HRA�K�W; ��ql�m����K��G
�Zy}ѵAF���L�2�5Y�p3/����
�(QB�z�����C�F��WO���6�e.��o�����kO6 ��*Q��4X��n;`M=���q^'�J��Mt�i1 ��2��R�>���Dj%ˮ��V�ȸ�Z꞉�C�����gڍ��-T�+�m�ѝ9�rD�ɑ�W~�O�h��M�	u=��K�E�Hmr2	�{�A��k�����c�uT��Am7gW�$�t)��5��BA�ŖQo�(�>�5�M�'wA诋�oՑc�r W6��h��Vu݁DL�q�!|qw3Я�b��v�\��0ш�,%��pht��?���t�Ӿ�?*�*$�t�x>��������DQ�liXV��(��7%�FLr$���IBv�y���-53�k���|���I3��6��?��Z��葞f2g���f�}G0��s����=ѥ���)�Iw;��.�=h�^P+��jG$46�C�U���}� �<S[��|Ѭ������90zr�@b�S�fZ�҉���)��P�L�1J}R���/[��.E���@ʙ�5�?F�?-��5.��_���k��_���9V
�.C<A��<7��3 q���_M1T
�S��'T��P�-5���2�{��2y�B�Y c>�d���u�&ڼ�s�`�ܸx!������*Qi�����BY�� P�8�:'��qi���E$|�3�#���ָP"%�CJ!��R�"M.� ��洂:MǐF1O.�,��Y��l���>3N
�nؔ�l����]ۖdW�:7������Q7Ǹ۵g�MhRq���m4,�#tE�9���ǟS
|)��F��Z4�(���%��P�)k�ZZ�ф�����R^E�!�ߧ�́3��BV�k�B"�#��M,q�<��dU���)��S�WMr ����~�Ѳ0�Zv5����b?�o�$U�VnI�N����Q�zU̯o���꺳%V���:����[mb �<���\�'�&H<?�x`#�؜O5\��1Z�&���̡f��m한��	!�FYV�>��c�e�ol&i�x�|�,��A�Bo:)�?���6J�
��ҼV,�LT�d�S�G�XC�*�!����M�C�D͜�M U�(�����mF����I�J��?#,P�؜45�iFK��U�_�(>���Ѳ�%�G;��2W��n1q�2S[X�*�����o���!��C�ލ�>8�ڡ��i}{é4NIa���sfJu6c����U��z���a;�Z���ļ��k I۷�3{-|߫׏����~L>�r���Ä�C��9�(��E�q ��G�v"��l��xs.����Ǖ���zv0���;�/�^e�Ҏ�Ҧ�Y1g~UB�O��ՙ,V_�N�T����E�=i�����,��K|�u�6N\_��"nU��5�KF��14�c�Gt�\��O#�vdB԰z�f��˗�����A���$��'��AC�R�'v�Y�+�q�
�gd�$���t��K�I�������sK�h"���	��%W��0�K.�|�xAX"����V�٦8��:r#Mܹ����¦�J
k�j��-�H4���6��=�/�ǈb��o��'���3���7�@���O8���x�OFbr9.�Ř�$�{��)���R��Eͷ�0�h��YΦ͊�C.��HV�]��)�ɷ����j��+-�(�MR���G�p&��3����1[��J���!��1��k���\k&2�w7�~o���~[����q��n���������W��Y�'$�W� '١O����>���7n�qB�tgt���"�CNn^W;�)���_�l:�R��:K�l�N@�5(x3�c:6`\N���S�M����y 9�pnE��*.W�Q
�����������bu@gV/v9��ۗ~�1X��p��)>s!���M^�L�D��쾄��/�m1&��MEM�R^�O]� �"�����}5h�~�0H����F#Ԥ{q��O*�)b��1�"�DA#����S��0��V�O����ÏX�s��	�!�KLX���mI�$�X�S�i͠qe�A5�@�|�a:y3���uONZ�B���ו�Ap�j�ձt0z'�FU^h1�,�}g�PjDļ���s���z���ag�+邌�o�+m��H��$����Pm͖�\h�M�-�4����3� c�m��!g�=Rh�s5�\�f�S|���D0��
�+uo�ɆVe~�\Em2��+��:Ƃ)j飰��6YO�����x��C�º���s*?>�"5ި6�����債�p"f��!���6J��ȸ������0��*eE� @ԦP�h멘r]+���'�.A3�m҇�� �W���Yv�TAz��RS���좍�Z�z���P���2�G�<�]�K�b���2!'0��aV�2���	�k#0���O���}P3���ǋ��s%�kM�b� a�8mL�V��ĉdۑ���]PKr�rŦ���)�`Z��]X�����e��.��v�;�+��.��L��?����d/������b�8�`����'!��p�v+3�n�|c�b��i�e�H��ٓD��E4�5�ģ��.��Ɗ5�H���S�c~�o�:;��a�Oh)�
���&�S`��d�G�?��F�������Gm�������'���O/�Z���t��-�iy���cJ�*��N=~g��q{LF���DA�n�������_�
�6
�6]�֩�t�R��K�?���M����������lm������΀1�(L����^\��w��㡺%W\��.s�<�����ܚ	H:�Y��`_q���~�������i��HM�s��Zop�g�I����خ���sSG �<�LD!��z�Z\L��P��1�qU���/���?��6�g�ӡ�����������fa�����&� \[�߽���x<��L�,��>ɡA͒k# ������B�][��h�Nu0�[A�H;x���R:�\5�K��Ü�z4�W	EǙ�*�yF�ݣ��~߼��,:��_5+���g$�i�Ebs�[�S����23�穡��z��1f��8�{���d�����H��ỳ`t1I�Q�Y=��=(j7F�: .�*R"o�.�/m]�[���Nuh������X,;��� C��'nQ\����P�nJ��`mH�*j��^��� ���LL�q�dc�޶ơ4c�#�g�w����%�HHH��'�s�EfUp���`�{���홨TS�4aY��8�q�	�W�脒�5�JP�8�8LS�Ï�Я�MQ<��Q�@�o��[tN~�"3�S��f��cj�g�� D�>��������֟L�hK�=�	�2�9�_�ʅ#���q,C��M*��J=�w(	ǟeLH�I��^%�\OԸ��!��P:�+�v�c��j�29ИZ̾m��8���a��ؠZ��~\N�cw'u���C�|�y����	����>�_�}Wjc�O�}9���愉6'�8�����N{�|[��n��%߈�������c;s�����xg����C�bg[W�$�w�%�{b�E\���G$�)v��TXh�W�7]��A��	'Yn���Di�mt�"�2s���P �e��_��q��/�WB�5%��0�L��5��!�j����?�XL�&�8� �CZ����'�sl0�ڭՌ�j_�Uꯆ��X!+��8%S��I���	d�^U���y�	��$���p���a��<ᇴX�������<F�j�z��6�-�5��u%�b�|�g.3F�[�z��?\o�x��:[��d��g�\�'n8��Jh��;��U�����iFD��/K̽QÛ���
.d����!;Nt?ԑ���Rۢ`�"33�����j~X�̝�qy	4��KS�th���)���\d�DԀL���y	��;S��l��k���F�}��oY��˧(�y��@�o4TR�7)=�D�l kv�F�%<3U@T؅5��t7	�G���$��k�ڛՓ�QͿ��?-B��O�a�/}:g<	�	ЍɅI-�TF����'ء>(hy�[�!m#�(n���i<Xu��Ƒ�@RbA��P���RĔBP����s{��|�x���n�M-�������|V%�Y���k�fȖ�����]c(��-��� �j��I�@L��ٿ�~^A��gI��3?�)(�Y@���#|�F���+P4{����c'�R�����~�1Z�Ʒ✟A�����|G���{�r61ߺ"��|�Vƨ����&;�P$�����9�+tji��#�b�`��縒Ȝ�2*R�nY��n�k�7œ�z�!Z�͒(n�����o;�6��ʳ�NA�O�-�ho�&��-H���7}��~�׹�P��p�ߙ��s3Y���{0>A.|�B����wv�BՆK�V�K��W)*��j,	0��x/`r�/?S�6f��<+���=�3�y8Ѕ��{ In�.�V�� �4��͔1]X�"Q��,�%�.��t�ov���2��g�X�����<a��𹙑E���������l���I�6F���B�6�|��圥���Hޯ>��E��FҕA����t�躠Y
��L٣]��q#,���V���m�����B��ҍ��1.]"�Xwۭ1��qa�;��~�]�qW� X�+��vRT�fG�?��g��P����e��|uM$���K$D	��&:9�1����A�WT"��;K�3�nn�St�և�f�-�a�4��	��i����^�I���L���"A�T~9���/��	_Zx,�3Y��rzk��
��1�.��b�0�O�]�h7�s��a\<Q�i/���O�i�������wyBb��!��c�a�f��'UfLw5�ҿ��puPmƸ���2�m�C'�ӻ�L�Vd���g����t����Pl���u}��8��$]��z��C�2)��栈���s�-�I.�O��i�sm�"6w��Ă5}[���e�9�!,��j���!�o|��9��ʆ!�����z)p�aKh��$?'��YJ��;�"�u�kvn%����IeDEK�"g�>N*�V��O���;А�x�^:�e�L(�!&��Q��<����Q�_<��7H�Vc��=�Wn
���� g�p�3C��Z�o~\��w<rF�r��ԍX�Bk[Y?���t,='?C[/��c���y�E�u`��a)��ل#`1�H�H���|�A��۰z���Y�+>�`�A���б�E�8�w�.�|�3�g_ٺP��P	PB5�&��%�dB��hs"Q6nW\h:k����sp��'t��&y�aDAh�Z;O�L�]�jz,,;���F!�2~M�2�v��ł�����G=S��u�	���6���W���Y�^��`I�K�&- ���d��`�y�4E��Ѵ�?�� \�E2��G'�y8Đ-s�ֈrQ$�༫��:��K�I���L�Yhh)X��iqg�^�?��<�L�I����� !��G�ܦ�ی������������N�'CѼz�Y�I�`7ʍ�0@�*6@�M��ߒ<�z�m�3�9A&�f~�	n)�H��S��#�]�������f"��N-��/1#��'n
nR�+��|Ͷ��١a~��	@J' �!���E�R�¢=���nR������tP����q#���zX�۬���`ֈ�MŇ�[�l�@�I:p[�sF�����Ϭ7m*�Bb"6���l��߬j�a��[���Ũ��㡻�>�x���XM㜁ۜ�O��X��A�b�L/@��\l��}�����{qI9��o�Z��i7I�CkF-?^��ݽ[��_?��x�����y����^1񞶞w�(M(/��E߂���%� %1�Q���0R齟n�D3{%�U��7���$�������-�]u�B����_t�]U�w�y���~f$�=�Y�|R��C���*hJJgc^J������נ���n_ hD��S���_�a�[<]XPO�YJ���þ,Mɒ�D�W2�Z�cD.�ޖк�sG �
�*tȾ�L'��uWI=�S
�o2�)�k�DA{묔�&�C˶^���*�)ҡ���=n�:�B���&���h�ߺ��O��U�$�����I��|��d�.1���=�..�u�p
�mB���.�w�t	���F���2�a���wce�pF4;'��EDU���ܲS����-Ѹ7�/frX*�k�&���ү��7�DJ���4T���N	�G�	ܗ*��$I/���a�uaΔn'c-��|;�$��g6[M�N�%�z����2+�g3'�bg��� M�oG|��5����r���%�Fy�-=��'E�C \Ȭ]�V`���h�"M�1<��=�TӹM�7𰥑��݇�׃GUj��ΞzF��]9D$ Q������t��Vh%�f�ZvG�iY��W���eUbm)�K�ga�u	�V_��ڼ/�r�?(�Uq�������M������&��.�� [qZ;��z�zv}�*Eh|�}#ww��os�Ð[�J��W�Fv����%�&/`-s#k�rVE&��^k,���@��m4����=������F$�'3�e��e|�,���;����P�=r��0��������/��ʁ>$��Δg�)L(���i#�X9eg%��HO8f�A��a1�z���?�t����������v)A�������Â�٠9]���7�SfE�X�m#�x/P���@�����g�����W��v�%I_�?��"�H�W��b�h(�t��}w���*��y������w��g�:U�A����c;��c�@�J�F<���a荥�bT���>��Ҙ�}6ȳ��_-s.�/0��Nq̒1�"���q�yG
��J.4_*E��~�k�v�R����@���F�b�̓�@�c��^�d�q
ۏE2L�ҩ�p�b5��Rs� ���ٞ��H�I����ܗQS\���S_[��L��R��F"u��a�@^-΄]�F�����{Q�������	��S���]J�Kt���5���ᕩ�M׊^�1�,���@�X�����{a+��E8%y�MD����$v	!d��`.�6.*a��2�fAO�һRǤ��Zd�^8|Y���ٮ�}7L�)F@�^�~�$.6ΞУ��ՆP�8�H�ݹ��!oA�q���?k5,�OP|be�G� Ѳ�h������kmt���Ɗ8��=���8��Wi)�������̗4�{޸�7F�E����I[x83����]����/+c@+�熲f�����>��,���m�?Z��,P��-d�L]��u3;�DW�_�%��2g��Q62;J�nbA�r�����M�eSm9�#�)s�Xn�mdL�W%k��虰�
�ȼ�-D;�����T@��޺��zp2W�9�A�:>ŇXۖ��2����6�.���k,��1��c)����$"���� k�:n1�L����i���(i��L��$Ԋ $���(w���:����ĕ��0��hE�*���$��:��^R4���T�`<�'�Um�6���ݎ��2�}I(�s������i���+R
�;���c1�ר%c�>��O���[�(s۷�Sb�ab��y��X�>S]�޽��(��*����yc-�ֆҀ��W�`Z�{.x���2XX��� ���+Q��!4���S��n�_ ��u��^t�1��X6u��T@f�����T���#�K�>a��l��Mǧߡ��	�0�<?�z�W%��t��gEF&�n�u5Sl��n���В��Jv��� LO�=d[�U�¬�����e���Tu�>ӏ��n�O���4%��C�aO3�u���^%ρ y�o?A�&�Vf��q&��iV�x�P�7Lz���"�Z���&!�ޝFM�W�Yx#�܊Ӆ @w�?��'*������V�����	ު6Y���J�9a�����O�	NXAb�%?[���<h������Z�L�0� �E#'��wx�g�O��{dB���^�^0�NP�,7�b�R{�N�4����f��p��3=W��HHI�7a�t��A
��@��nu7H1M!}����IQ2OZ�8K���4o�ۢ������/�j&�]
���hRd�KY�l�Ů�C�� �s4h