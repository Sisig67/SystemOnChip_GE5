��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��׶8۞�@�\ږwiܕÜ��=r(ro�fC�pr�L�O�q�;��?���d��eZA� �t-��-R�l90*������N����
8�W���(�q���2��#x+�nt�,m�=ῠ���WDt����Vӡ�]��Y7�Y�6ڽ_�`/"K�X5C�\�h��tA	V�C
 LY��ۻ/�UM��+����Wռ�q�>`�T^��@'ʹ�H��f�h��X ���S�����#��n��hNg�}�Ȃ�s[��KЬ�
r/�lG+_ϋ9^ �Ɖ����,ެn�e�EY-�|W;��ù���=�5���mA�`��yTj�:~h�����#��Z����Nnu u��U�,����a.�>�1�������68�厽j�ޯ�'4v"�o�I:�/2I(�h	0��-�AW	��%*���Qc����1��3	���.�ʥ�rp���'U��#T+�&�73��$���s� ����xJeS�)o���@�^��C_ӊ��?�3긋��i�����:��w`㖲W �}ϼ �
uZ�x$�ko�YI�QBx��ر��Q�y^��Ib������v�oc:`��N%�3����!/�ԢDj�x|�=�� y�,hy�?�Z�f�\����X�V���]�N���#MVҠ�0�Ev����R�Ʌ���4i�!>��c���������Ƨ�/㝹�r������x���t��#Mp�{8����qQu���y"<�ގ&���q������<?���p
<�5�4)�iC��x9�.�׋�5��8s̃w 4�?vpw��ЩT�a�1���e���WY��d�M��6&M��'B�17:%^�8���4](K#$q�kȋ5��K�CO��fB������:ۄD�;������J�Sv�+�����[Z�_����b`�i֊f�{��f�3�=1ؿ$R�B���u�T2���_��݄�1�̷\ ~?��ϡR�]��8��Z	��C�9�)uP[*���d1
b��}�D�"��zi����o�G���0�\3>|Վ�E�c��.�3aYh�=خ�g%!�;�cE4�:>�{Q�����+& :�����`�,��k�������~�Ih�z?�z��ǁ�3�6��y(~!.� �Bw��o9%�6$�HԺT��e�b���?9ZEJ���Ͻ9���`
���ֈ�dgiJ��3��%J���xϩ+rV�n�^���͆���)~1����!�sg�rY��8�������>��5�GL�h�'��zɴ뿓r�[�i#,��5zH7}�G$*_��g�4�&ek�OZP!���9�����ݛ�_+^`��^l_�$�b8
���y�U.�I9��.�ESܖ+.s�2�7 70E�Fǆ�� ����$"1�to,�@��s���<�/�a�"���@䆋��/ց1��!\��Y._��~��UCD�*O��$H�Ƭ����Β����J�] �[���IzlG9o���Q�&�����Ð_�1)ȇ�k{e���[�<'$�iB�"�������������W����͖Uoj�vmւ�y���|Z+��^�bX꺳'Kǝ�|��g�[$�o�����Qu��37gv�<��z`4n���i�1c������C�߬�k��C�e��>��*$����wX��tW-2k�o����gCX��?������w}x�xOr#�T/wT �j�{�g�I���{��v�k5�����k�e��s��"EL ���Z��[�/��8�����4����� I�#�L!?�[��:>� ��-��+�X����">�ft�-8$4��U(M�9|����U��l�E�W#,��Wm�{̰z���G�%��dl��I2iBZ���J��-TӤ`/)�Xj��/$�׹�B��ӥnU��^�&~�O����Tg}����>��uBܪ4�t1�]�d��Q��yW�
;xFC9
c�(�$j��^�;��;f��b�O�gA>���3��ߕ�%=C�7x�o�r�s)����L#D��%��^�b�k���E�`�8��:<
6��������z�v�n�ϴΐ�w��8��BW��UB�0�Pܸ�
��Uu�)u5�/;�CL��c�ո�����H��>x�3��+y��F������=�?�vX/6:@=Q��}r��(ĉ� Hʊ�?��#eG�����O*��oN�d�/�%áZB����^����7^����P/�yܚ�m�]��$��.�_-��`13��!�����ԧ^cp�(�[	}���Ei )�,�T&�w��Kg��Ю���>P9��n"�K"fl�۷�+#;B����OF�*s�����!�x�p�?���.��.ļ��\lРUu�鉾N�WUW)A&Ԇ�6t�h��H
B��=`y������o1~�P�4�=��ı�\���)M\�-�$�f��!��	̢I� ���>�}Y�>A|���h���5�HW&�	p���
-����M�^Ω�71����8�ȴ��1�C_���ݙ{���
yZ,�,	�Kt8��>V�8|-@�r%-<�|ԛ�	��.< _;&o����7�c��Wx�A��x�m�e��j�n��S�ٵtUn�Z���6�	��B���1�9�J��j�K�k���PwcЭ���7��X���9��1 ����� �\���5���NwŴ�1��Ư���7W�^��s����=�n{�8(2[�u�ᄽ'ہ�7h *baƌ����\ �q ��2pn�[/ȼ�%��*��$6kP|��j76[�>��ej���1T[�IrJ���]���C�;��9�����{�=6���<����d�(T ؗ��.���!��ˆ����
�k�"���.� ��n ��3Iƴtpv��W��'e%z�tlcO���DA��t�e�a됑Шz�~C�O6 �����F'�p��t&��$�$���F�:��Y3�BD���cD_&��8�KAb��cc �I��M�D2�E��?Bg]�es�R�$�bk��]���ĂmP���4n��-(��Ոd������\1Kx��ux%�
8|ix��ʣ�a��`Nk���{�'��Q���;�] ��v�'��=�&!�{�l�l�A�m�L�.Z�{:m��Z.���J���f��c���z�>�;R���"� �|j��?�@w�V16�6Ms�k
o*&��S�䩦�ʕyIY ��DV¢zl���Jy��Pb"�ѫ`3낄�U�"l�W4Vy�\�p�~G��2�?�|�ޟ����yYF���()#�c��C�Fuj����S��UK��9�T�c_xy����]3�|H��qh�=���q���jf&�u�?[Rj?���҈��}~�m���;��P�~l\/\GZ���~�*p��w���J���̀�0��R���]+��0��F�oN�M)&����_"��[��a5~��̮?�O,�㽼~�B�qn�v�'�&�$%�x ��G8|&��A\v!nP=�Tt �_[�b%�Bc���tڶ��� ���R�_� ����d�ǌ�&;���*���������,����ݼ	@�h��)n�6ޜ�H��h�c���M ��˺���%��*�u���pX��G0H�z����~N�j�����ň��8?��v�}�.�n�'󕹽��/�:9�~�EW��h�in0Z����~}��	.e�+�'�Er�[��k%����Ę�;"\�Ϥ�f��I�xc�ɒ&���V����O�qs�[\��;Il`hF�e0��mz��]@�0�Z����ZEJ���6��\�y��V]�/%W��o��Pfw���Q�W+���N�]@#������ኗ	�ʞ���YP��[�Es�*�͓���J������OY�'a�1�G�,פ����ao��,��N��pYv�`��`�.i+9M^x��c+(��K۲L���'ӊ�_��(	�1Q����84�+���1#�d��+��������$��v�`��l���y��{�H�Km�X3����Y��|�n����t�f�K�-'�K�q[`iw"��y4*7������;٩�����Y�F��ff�`�Fـ�.���%�D�~W&�f5��v������K���;}�޵̡{�d����R�� ��ͨ<Z�{u��|���ԗ>�(:.X�����������nQʋ���b��
���dv�I�[N N�B?쐳��Ѹ}�F����9	P҄>��nz���C?�
���%�;�d��0{�6W�\^1ڙ�r���6P^��A�.�܄	q��P��?�I�k��jͪ�<_\����[�t���f�eA�?�"��&���,�/v2̉�������=��������H��<�©׭���֚k�K�Rv�QrS�Tc!6��E���p�EK�ӘKs H�J����ݖ[����u�S�	G�7QB���MY�y�X_ك�$E�8_��&�_���)E�����$+䩧<�,�9��2���d(a3�}��`z�K� �ܐ�
�(�;�y"6?q�VU����4+���+�NXu	b$Oc/O[������(��k�TeD̾�P�Ĥ��vv-��� �fVs���[�<a��Ԏr�|<���G�O@�r����+2�"��`ݺ��%��d�"��5W��m7$�鶜�����e�Xmq;c�����E��n�� �q�h�R�rO�dG�Ͱ[u,�і՝Aqw�R���¥��=�q�+<!V���i4��Y��0��)�e(���FR��fPe�_����j�p�'N����gӐ�>�����Jg��ZDϵ�l`�`��H{T<�*A޲�<X=G!���۞� ��H���s)"�V�1���Y�I) m��$�EV�H�Tm$O8�#`ו>�&�!��w�!��q�2�����*��$,p���������ɏŒ�� �''�^��05,����Y����Kğ��b�ff$�����J7A�"�� ?��xm���y' ғ��&cN�� ��;,]\.�c��C#4Y����o���́���-�EK�^et�}h����V��]���m���7+�9����˕K�^�v)�O�~��S��I�'������p�$��p���2�$7�ɏ�\3@��#��~�8|�B�~� QqͰ8�,��ڷ������p
h�#��/}�W�V��T���B��s���Tb��I�U㐎��V�@��%ӻA'�4q^�.%Yz��F��:e��7M]�y��Ņ0lD��~a� 7�𲈜��#v���a&�t������ɶ Ը�(���ph�f�yނ$�?#z����Q�"���u�
nĆ�7��'$�~C�_��i�b��z�lm`��o���pZEH�P���C��E�p��(����4j����[����i��bs'2'ɼp�#sFF0^!�rƖc�\O������xu�O�j�G�5�d�uLW��RJi���j���X��ke=Oѥo�Z��U��FB|�u�%��e�R+�Bԁ��>7g�h]^��L�\wTK
��Bz�W�U���!k4�t�N���{�Ͳ�d�l�B��A�\g(�2�O���9�+*�� �O��-�u=����ҏ�{@���Ӄ���S���j�)�J5�H�8ک��x�cK��f#��
?w�%��"�agT�J0�R#6�Ȗ �5{qΨ6�R�S�O��m�M�)�ع����C�W��Ӆ$�T���p\�Zµ��8�R��b������lf� �L�He�#����Ӆr� ь�nv�Uu��a��Y�'?qH�9v|\��x_���X�x�E��W��<*��B1^�ݼ6���:�2\� cd�x���_L�H��?U/�TAo���o�%c����6ӠXj�T��W�AX���б��Ju��{�9�#�-�;�=
�x��7sD8jgT.(�Yh��m�g���p3��Z���Y����K|����O���	��v�`E�
\%���^qGs�{�U>��r ��Z�ge�6���c�k[������������n��D<�'��ڨ3,Xh�yV	�*\�7�^¼|�<�SH8��|�[5*�/Nı�� �y`Ŀ	�+z��b৒Y��A�K5��V�=/�"�=�'��9����(�.9d�@�[�T�H����\���:�jQ�/2R~���FS�Y!
*���c֮�x��zLT�1�VY���DQ
MM�O�&u,B�7�h����2��t!��t���.oZ_�</!倕���u@�2�'��5Dy>��"�S[垺+|���^��iM'@�2}����1ـ�D��ĕ�9������޾���y0_p�P�9�������7����s��I� )eCP��&���@�̫va��3+�l���L ��q�g��@�P;%Z�������*�3��6f�R-�8�wn5CN�s�˒��iO����13Ar�	C�r8�aRu=��/{���K�oJ̸���2y�X��]�����}#�:�[��8���iD���L�9��jP�S�f0g�)r�W���m�X"u`�|��<H	^�(9�4�i�d���<�G@!���v߯�l�^�*���o
��4�/�}��M�`%�J��A���#�B�?�r屪��7>[���w_�:����T�yq�7qk�	]��1�E���=ڣ8�� ^]o�3�����r��|����E�&���7��:�y�Rp�.�H���G�3�9{&T�jM�n�lk�
i������e����"\҅�va'��3gO �����>�j� �o�t�4�+3��h��wHZ�U+�����\����̇=��G����3�M0h�J*E|�} ��e$�^�
Ơ~�ʝ,�����!n��
窇A#�J�?!� 1�Xmwj�`���?nz��$�C��?���fRc���d�E�;	�����UT/0)IOuH�ŤƖ�2z1� �P�d���n��9%+��r\����N;��yQ��u�@����lo�P��������K�9�5�`�����t�_d��J�q�-��`�z��>a5?���d`|�)F|�7��,�>�ƣzL]qĖ08͐;bD�D��L,�������j�,a?L�%���>�{�Y�R/э�wY|��dCM/�4���w�۳�������
z�+���0��\Qp��%�^��IR�d�#���9J�t���r̨�����S�BѠ:\^�_r�	�}��+�==�����j��m vȆhQ��ݮͤS�֯i�o�(j�w��j����;=e}��5�E��OWoUy������� AnYR�o�a��Q��ʓ��A�O5�y)���!�@O��wq��J�{��H���йJ��$�Q�����Оg��ٔa*F���F#��1?d�q�²,�U�- -��a��t�OIR��qo���λ��5�'I���)�av��������Ч��QA"`�	2S?��4���Op�aX��=/wbC��e�,K�:?�r�0Q�r\<�k�Zͽه��X�]��g��L���b�'ؗ�H�s��N�R`�>uX�K(��#��D�����zj�s����l�;v"8�5{Gq~�i��R�%��%�Zq����d�W aSm4Q-W(=���:�&�䍚����32\0��bF
;�`����Gt�o���3�qI�G���]��=�@��"5�vFTmN%x�E*���n��52_���h��u���8B5�-��Q�TB2�54;o�M�	���ꕢ��N�?Ύf;�k������D>�N�bƸ{�g��Sq.ݧ��$�춟�pH!�W����6I/��>o��`Iy�	Rd,��8,���K�ä4�bQ�<Qk䜤j�~0?�
vw ��z/`\�O��x��&�X�B�~я�d�����a�����ס`��ȓ8Y�:jl���A��շ���/���yo�����Q=w�a���k�	�t��PWqT\1őE ��8�"1냔�o�wn�{pi6i3���=jbb��8�<s�i�e�u>}Jl��ς��%�J~]�bm����h3����?$ÏJ���<���n:p�K�W�<���d�ˬ{J ����k!���8� 9Ѓ=�ySZ��4�Wc*�K
�J �O��W�i*[�8K�2e�-�gz���(�/h}��� C�&��){|4(�����|LN�{ ?��&M#��Q;'z�4_K���˼#v�_�K��W�ʪR_8�䝟P	Fb ������q������/ѐ���Q�*���1��C�"V�B37O쏆C��>������L�~�όF�P�a�H܁�r(�q��x骼'l'Ţ�(iR��{|�cA�O �,��w�ZΩܛ�08}���#i�8n�G�T�D`,����?��|��AH�J�W�[���ωA.�U�6�w��6p�Js�֋K�8"B=X��]�P�X��0H]��6�T%ڹ����(�{[��PM�τ?����;c:�����I"�ց�u/���)`�K#��A�L��v���~r���Y���ǵ�!�����e�%�_84�"��j��1uY۟}g!������<l촰*K�`��՟Lc��{��~{��kVdI���i� �K1�h~#�V�ݧl)�M;������g�z�/Tk���7���{`W����WV�4��gR\�!��`��ہ���1X����ͥl�"/�n���)�ٌ_������>��ob =�%�+�a�;��ܩi�)�/�~���a�XUw�N���QH�f�e��i�:l���y]�7�_��\uґ�-.[Vr�
�����7T����~dx��a+�����h)*m}1���V[��5�����#L=q�䢽�(�bGZ�9�� x�TV�K�a.�^Q�1��4�mE��gm!'�O�H�K���K��-���Ȉ�˼��M�y.Sx��f�㗊i��;��0�t���/�:��M
���gV�ú,q�ٸ��ނ7���e�a�� h)�	n`�����
��V,�mè�Π���/Trk�HDZ�o����W�o�����,����	c� �� ����_�,��ǈ�E��h��v��QuU�J"v�:����Q��	�t�.i�P@�3!��ަ\ȿ��C*�紷��m��4��l�6R*\z��X��P��$��3Kw-���T������쀆R��Z�G�F�	> ���I}�#�er\���y�a2R������6G�z17�$B��%������%j��>Os�7���
;jb���u]GC��K�M䨠۫9����vi�/���K,����CFqae���\>Wc)�@��L�֔�1L�b�~� ���|���N+��:�b����"QHz^G����dӁW�\d��u�Bt!D�Y�T-!ߺ�Ig�xQ^��b�&g(" i� Z�3�yP�@J���?�T|8{i��U�z���=?�g�H�^�3@���'��:�[@�Y�����8���6�ю�}l��ϰ	.��'�C��4��\���K�����.��+=eHZo+ �6/D��(���Q����>UE�<*R�N}6|H�!o���G�9�Y(Vz"��i�7z�O,o
�-r �$|(�S	�Db�pj=&���i��ٗ�o\�h$�����⁬��N�B����*m1ԫw�P�z�(@Zj->I�N5�'�~����Ė��E�	C,`���8���*��%��z����*+��ޔOM2��O�j�R<{,�)�_�[��j�:��HҒ kR"Ƅ�v�Ld��?%��`��0f�]%�|q��Z��a%�u�zvu�K��$~ݝ�H�ǜ����z��5(���,>�����b�2*�"\� �����Lu]M����!l1ߘ����J�����ᥙK�������}�̢�����m`T�T�Ñ�}kb1�Vj��9[:�0:uT��)���F�P�V���x�)B!�i�iW�4�*�5��ø�yU��~s�N������l����P�ç��H(�N�Z[S3mz���A�E/���^'� ���aँ�B�	�.`G{��&�h3IX�#�����}��C��~�u��G~��gt�@������TZ�*J�!j+S)P�_U� ���=Q,�I.NzmS��q��^qAP.@��c]�����lP���05W�L����ct�Kˇ$�3��K�Y��Z.<�ծԎ��l�b*��(�<8'�j�� �CM�^���YU�zy`�����uS�e�s�w�G�����I$ٓ�Вsq��c��rMq�NTZ�<�r��F� �c�<=���Ğ��RT�3����1�m;x7�����>���Xj�Հ��T?�^�k�޽j(gܤ9�XT��
��"�^����"5usm�n�fpJ������@��6�;Z�@��]�fO�B}��\�&�S�b�i��L�a�Z��(b_06��Ezu[ӳ�� p[�!�u�&�&�g4�#��8:!+�-�m� �T}5V���򜥑Q���e��׷o�!`w�w�e��=k��ԊYBz2�������A�%~�y@[SQ#8Y��f�+�
�w��hi��J�T��U�{����T�tOЕ����T,qd*'=IS��8tI�~�,�N`��3��=�m���[,Cq[����RB�~Ā�����c����z����G��(�bfu>��oE�GKc��cdoK�]�{ �NPm':�j&io��-��
c��`���5k
��wQ>fi�˫cw�})/�8�z�E����7�5�/��e��n����d����Q���\TA@�z��6f��F����nx5e;ҩJͬp�P� ('�#������o"�u�e?�j߯���V��NV\�=��L�֟���i�R'�&3����i�LM���q='��j�'�|?`�el߃W�;3�Y�~���+��Ɔ,��Y 繓��y0�{�!w�-���Ў[�<��V�����N9���;\z�O���(��3�y}�7j��m�Aϓ��@��
xiqj7fQ�����X�pZ��l�[e}{%t��뾳+��Ƙ!�Lk�q3j��ǬLx垴,�B�;����P���Q?���2תEvy*Ǐ*۱���0s��Ǆ����Q&\ZƖ�b��Rx,�����l�u��Dɲ��9�7���ޕf$
X�#x�x�p�B+%T�+D^e5e^���/�LX�(��}8�L�~Wu��c����KPzݘ�c{�88�6n|���@vQ�$wVߝ��p��o�γO���0��c,��]u%�1^t����E�[h�J*s������ �p��+����<�KU�i��ݛ �ש��_�Pv"��XKo��$x�=�{%�Cl^�Z���?��d�%v��Z�Z	}j���-�kC��/m�Lh`�K�q��K>�T�E_rk�|Oڒ�(�����Ht1���j�0����l�0&�2��@���M2М��EL�T�{��2JU����6���+WS*^X`�Q(Z5�u��#�>PuTҟ��Jp�3��_�8�X�Qz��Dt��|�����%<�m�6{jC�֯֨���wr��]U8�F��S����Ѐ%)�����@�J��<z,��
Q�����k녦��ߎPju�6qq���)[�;0-�	/
�l�猘GU�v���
C�Ȉ˵�0mJ�ҚrH�u6�U����C8p䄣o�����&
Ъ������c�J}�70�##�kӗ��?�ڬI�M�ȻD5�T����BJ�`�s��N��J"U���:�m��%NN{O����"Oz.��]8˕#-�дv^`VdKŌ���N2	��cvC�t�[s���l�h^���D�81ހ�������fxM�O���OP���2j��>�r>`�vw4�Rڧ�a}&g��	-��U�� ����� �j<�4�-�hM}���=��.�"Z>Q\_���.��q/���B�]��T��?"�};���TV�}�#��ZJ��/HfW��sK�+��\1�FL���ȘW=f�mYe��^RT��,��dOP!%�y�/ݺ�C����.����yA�� `�ڪ��>�m,�0���o閺�a��|��=�EX��b
���ؤ�_d�o�g���u�0-�Nw�f}#�VI1��c~ɴ��/��Z�>Q,c��g0���ZGj��zz���e�!�qN�o�=qFM�g���i�,n�%�t�?m_ؚh������[�A�I�)�nk\u\�k6��,�^t=6>Ѣ�×�H.���8;O����\�ֻq}ϝ�()�N���k
�B'U��A�S�x�y�B�A�_aE���T�U����#��G��܏GK�L;nӏ�^D̶C���{�lK*���;�!J�X��vM�͝*'`��t�XU!�t��,�L�J�=n.������F�T��T��ӝ��e���O���3_�,f��'8��-F4%�`$��7�����J���[G��0���k�b&�'����5Qk��3v�;bl�e�m��=O���{���iC��<a�,��q�춑j�Ug.1N|IC�����4��|��}ˈ/�ȥ��e�(�	)=*��ϥ3��CB(Y%�wM��_�#G���ɀ��[�5���K�<Gg����FDY���F4����}0��t*��������]N��HN��Q�H{�c0-�
��_�����Y4�ݒ�0�S>ԟ��K�/�ȊDg�$��Z��{F��v�ǆ}Ygo�˻�D�q���ٸp踜�8-F��7��:4�QǼ�h�ϝ����o!9�"om�x� ]�e�Ã<#V2��d���>��g�(���RV.��EA�	D������Y��n���KvU�n��� F�%�0�+�C��ԢƐ��Dv��r&+�9�.wuG�6�G�NP�[Hs�8�u������3�[��Q�Z#��f�)��P<�,gN���g/1�&�4H����$��8�{key��|�^ѯqC���gD��J퀫�xx���R�h�a�N�ȸ� ��R@R���^�FC�j���`���i�hUL�����x]�|���s�V�,B��爋�]���yYx�N�>|e=�ߏ���>�N�L{��h�q����p��	4�ކʰ	Pd�"�bPIasz�����F>膝̀�;��N�ks6��+jףּ�W=XD?\c,�]�ZN�f���؁��0��U�nK��1���2SQN/ W7��;H^!{�������_)&A����;�[��u�P�BGRCK����q�叙u5 m�!�+Ê���-��N�_���#�?߇7䮱�i�� e�Q�FOc�8��Z���~#�,�f�2dڈ��I�evދ[��1��Gr�od�JԞ�w�|f��IZ���66,�����P�>͈f#N7 qP���D��t��m�m�~Tkwj ��qPT*�{Wt��$#=�染�й5�)���5�Ɲ�R0���������BI�����k2�a0�as�y{��$��Ղ�
�Px�j
۲NjO������x�\�ԗ~� ).����SBuq�-ǔQ��ҫ9���ZMϦ4L����
v�`72�%Rr%��#pQ���u��������+O�sʟ���BNCFl)e��N>-�
y�2���	�����
;� 8T�	�H�%O��0��
N��Z�d���ݚ��:���|-�y_%5Nk1��*m������|�$<�\������E�09z��0SdN��2���c��fd��!������^�7R\�y�*�J�|���86x�P�i���!�ʾ��ZUZ#c�f.�7��	
%m&IP����K1F�4<���J'zD<�TVai�5���z<V��S����<�7m��1:Qv�@m�ȝ�z ۇe%�E���b�~i!Ui�"�$���L�x�����VI�a�^A@�3L.����p�VĘg���D"�]��A���ɿ����U��(����]ܐ!mc
ߙ�i$��R>��5�3Ґ#���)��s���'�����\�}mִ>�;�r���=-{�>�����C��[��"�
7��8�25��YP
ŬA�򥔹H~w�3��m*���f���n�Z���d6����q�cn<u�f]���^��p~Ȋ>��R)_F�,؈�:m?c�������
��T=P
X���O����� ~֧7)5����r���k�/�aYۨ��x M]�'�/��MtY�ӆy�*O/{�k��sHhxz�63g����.�Ϭ��dBG�]�����i�W�
�ʗ�ɭ��j>iL�1̢˺"{�1k����*�y�c����	>k߃�jgj��]�-�]"�]�b^}��������pC��Oa7��c�(�͙O�2��i'�3��2��h���1b�	��`�A`������S>g �Иƶy�F�2�➧�EE72�'ؽ�練���T#��׵ '&�`��[MG�Sف�o�V����aP��e�����B�yP�6�e��xn�.�˯������+��|���6v��[����t�o��}x\��ϣ��
/�v�̚!�̲_�BEsv}��J���rJ@^b�Y� lf|�m�˿!q>��)ج��5jzÔJz���j-b5�Wه6V��#�%���LP|@	Dv��^mu�ϧR��dh��vbWIÇ�$Ci�eq�))��q�遌�ہN��NSp)9�#�^�{��Q����b�Y@e���V�O_�-��n��8��o���6Ya.�b�I=_-v��HF�3�q����s���u:��,�F�_4��ze�q��JςXZ]l�(�[�y�v�cŊ�ɦ��iC~L�9�3�Z�qZģ[h�ui��p`��$dg&�U����L{0�)_N�E�yW�T�GN�o4�U8A�MX\���Ga��>���P|���3�\���e�?�F{ޜ�gW��1�L�@0AGR4Ф0͒U�j�9�W�$VF�R1A��Y|.���W`�����OQ �� �(L���$rv�&�`95��u���������	I�S�*9c�^`��3�,P����d�����*]��h,Y��c��*+�o��u�����h�,oY�8|�_L���\U�)Bq9.SV�t<�ml��%a���i�Q�ϔ$��N�Y��[�M��Ցm��sS�t^o�I�K��/���F����;F5�R��/�0��\�ѝ��o�*�&�@_[��8�lJ��;]�Q2#�C��z8���}ma�56z7˚�:\�F��E��;�����D��WT���WJ�ٶ����ߺo��?�F/Q��/T�D�4�������YA�ǳ?f;WDb�L�7�*N��?zj�y��B�w�
�"6�_a0�������]a�[7ˡX�H��M�+�mA>�7���0���p�&U7�~��E��a�Z2��|t$v;��]�|���Z0�h�?Z�^)+e��Qy��!�8j��2b��V�ʩ�W�_�A*��8�z���C�*�u_@�c�C����:��\O�6v�6���-U3Unt=T����x�����՘����^Ll�3/ꖱ+׷\ƿ�.�@*����O�=�f��`S�ϡ�Aa*-~茪߷"���+�C@����c!Qs��n���Az��Y@2r��FQ�6p�ݰ�~%u���X�3B�$z;`D��/�Z���������8�A�a�HG�X�r3k8��X8a�����D宒�>�y�wwTԫ]�w�ʶ��$��3{:�.ȑ8��[vYW�S�M����~jZ�9�k3��Ԍ����%���b���(�+~O�6&�a6Վ�kՒq\Y�%������	��[ꋷm��p�2F�j{#] [��u�1��O�A��#�?�)%��Q�'�J���F:Z�6$��Ā��� =Ί�uGh��w]�u����	�G}��.�';p�,L��Ј��'�����ӗ�gr�hxW��tT�t������5>��:aEJ�Ҽ���z�\�k�:3���<�ѯ}������T��.!���V_������~�.�Y��|�P�Mu5�1R�Ý�vI;�O�u�sn0^�.�YT�>��l�����C��e|x�����'8�R1u@ěiq���| T��re�#�ᨠ0!pzF�(���Uq{eG���B��}B	��u��@W{Աl98l�)w����UT�d�5?)u+&1rol�'ft����i�%zkaCnr��;ѠJ�Uy�[��&�����xv���r`�k�M�H�_l������qv ��o�R��㥶N��">w�ߖ�e��(M"�q:�ԁJ�L�n�.�jE�������c,W|��f���g���*v��ߊpeYA���T"�E��L�&�dKk�����O�*o~o>�*-�Œ��0:B,i�ްt��S��s`�-�G�G��`���rM �)��-D��5<͊{��K���������V��_8S6�[i3�A���J������ [�w���ysz� ��􈤂�sW���v{�h��TY��J��\E����������@ܧ.i�~x�F��$�-���,�4]����.�<�@}k��t���8��:���Z�,��D��grM���]w]�z� �����p�PL��^d���-�,{iYޝ��>o�����/�s<�1��kk�%џ���B'��=	��ȩ��ܸ)��b�J���)a�?�`��ujKP�*T����B�N�k��b�fz)�j��)�nf����&� Vg�`뮀0i�;��D��i��Z�b�?��=1'{��vv��_k���!�Ӂ��tEء��U0�N�u~9߫���1|�e��`�,~Q7����?��1�i���n8h���߷�=Fu����DVΓ_O0��;�`�8arK$��6K�HV��Wu@�M��㏠�-��� ^,'�
��۹N��u�E�!�Vsu	
9�inCt��?df`w�X}g`n}�|~ߜ����qQ�J���.�e����^���;/w��̜��pX�?�(�ǡ5��s/4%���% UrŘ`]
������R�������տ{?~/0w���8��Ǯ�-���/_�e�3�W12�oYu����x�x�d�;�'a��t��@�����"����*�\�[T[>S�I�����QO��X�Q�a,��Y2�Ա ��$h'��%����7�v�]F���
W�leֈ;�[R����W��ʒ�	�>�v�q]�3V^�־*���N˺�g�np).��r�rO�8񢀆��/a'�r=���i+�����M��I$
���gF#N9��Ԥ�hF�b�ݦ@���"��!�M�@5�\h6�V9���ۣ�o��=1�l�' v��b�=�������� t4E�9(�g��@Q$=����艳�����]�	4[�z���7xW��䓡��`�=}�0�0�Z�	X�K���F4=�M���C�m˩��Jw�M��n�V�c�{{Q0�~���:Uμ��d,U!��\�Z�����`�G�i�Yb�V�n�E����L��������G���KB���[����7�/���˿����t�r����rA����gN�u�T*&�M�6�g�e���ܣ�X*؛{�⻪IX��|���(�`@�Z��^_g�ѧ��@tevf�0���vy^�&"U�m��l��������)f����rZv�b&�IE/Q���<�?�Wa�}���ڟB��R�Ř���94�[��0�q`?���s���S�1�k5���
�/0�w�ˋr�[,9<>c	�~`4ߩ��QSb���;8�L�J�_�:r���Y�����*�a�LZ���y�"�Y�`��#�Y���<�B�e��ZD֥�U_8��]bJ+�H5��ʟV�ŦR�-����w�qx<,��=�{�"Q�n�Pc���O�<��^ �cD�I>�$؏l�0N�B�S�]���PO��:��Y�# �,��a��U�2�,���J=��w��Q��;1�4g�<AOv"�<�7�;�g(P�0�9��h�d��r�0]�u"��ų
Ɍ�Nx>��F'�	Jj�)����l��X�"��
���$������ш>�t�%T��0t죢 �B����=�gϹ�?�g�'턆��>���M�F�Uk����_Yl��棩qF�~��}�ݓ��A�~21�(C��c��*³�p
`���_⏨qZ����f��ٹ�MOײt& ���Y�l�[(j.���:�� `�`��	��2�PК֭#����"�a,+c���<$��ʧ�&��W ��ȉ|�+�g�:�� �D���ssf 0S��UͽJYD}�%�I��yH.�x����5�Suޫ��r4{z���T��A�)��o}3/���lT��.r*��`u�N�Q}Z��8�\����V �	� �eX�����%���k�c�*�%�ſ�[�U�VP�ij.�fmB��Nc(U�)���|07������XO��Ko&�eT��0�gf4�\}?=V]9b����u`�|�X�׿S�p���́��Ǜ�����5���7��Y�����3�6w@G�V��_:������M�Uԛm���;��ƞ�,[=wVE������4FN��+�P,j�XE�;��"�8�e�9>��tf�➆#D�cK4f�k[	kb�_ټ<�@/�i*�#��7t��yy4w���1q�3^\_�ß\l�)N�1�WUk\�Y�4SĻ�l������m`�5NC.�U*~�e�ro:~f�2>����ѻm���w��N� �5tV���]1D1�V����k�P�Ɏ�%|�#L^�;�X��m��D?�8Y�Pv�<�MЗ<j�<���l�0�E񳤑�!��R�e_e
ϗj�/��M�f�by��ΆS�o>�+����HG�#�%�wy�m�r�����x�=�V��P�#z�nL�����>b�t�B
��>Kȩ��n��H�[�2~��/��+T̠e�^�����c���9AG?�*]���im�g���W�׷ƻ������pm�_�B|���x�G�t?�$�'Ѽw�����a5k ��#{���<a����T��	��D3Q�^_1�6��޿X��Eɏ�=v�K�{gjհQʡK$Ķ�J��Uh7��>T.�H�Ih74$q�\��G����
K$ȇ�O_ꭨp������p6=�2zeÐ'�.�:�����M\ �E�/k,|�X���n�����7�n�ŗtB�������!�5������-FA�-��eѪ�?!*�J��-L��4�1I�0�����؅5���w5��/��]d��%Ua���W+Ug��l��[ٽR@�J6�9xyV��47�Y�/�a��KI�j�˵׽���&�{	15���Z��"=-�u��I}��{Obqx�=����'8�e߭BfO�⮸����� 	
�񆢞����&�i������\�~Y����'�8u:,���:f��oݠ4�=�wf],ƞ�h巃���['�L��}w�1^����}w�"��S͍r5�r�� n���Ԑu�������q>��o���8���y��˿ޝ��66��l�����"������6�Y�!6[-"��8�����oO���r��DyrL��U��?k˱�t��b���k0ð�z�1w^7vw�1�y�=���հ���}������8Ӹs��R���K=ݙ��iG�:�Z�Ȥ/Z�.M?\��9���
$�~���+AR/�������u$�LzP���RQ�6����������2J�3�[���j�ݣ_��!jt���Y���f����B>�Kҭ>�ܥ���4���+Le�P���O������1)��q^@73�.B����.�Ĥ�Z"�����~Xޥ�	����c tw�Q!���:K���!�H�Bŀ�Sx��U�-��8�b��se+�y�� [�i�9�&������B�`��y�z��F��j���J��uJx�0���ҧ"�P����c��GO�N�Xtm���9�b��g�����r���6Z�9���3!��������%�] n��7��-� ����N���ϊ��F�A�8�;��G����YS:�M�5� ��3T@�hy��
�OA�>%�C�����}u�EԸ �?���S$X������KL#yC��9���R;��UՎ�)��ʃO���'j��d=t§q�X눒��pqy˘}}��[7���%p� \�.��&�W��2��j[�D�_�3U@�E%�m.t�^��:+35ȓ�x�s��翄:�hv仃c5��2$���8;�.c�]�K���Ԭ���3P�m	�9�\��ǹ��/k�q����R.����	Ћ-���}���v,$�lpT��s�@]�ъs7��Xm�ݡZ�S���.}3g��? �$�J6����g�X�ؘR��Z��=g�}C�-���Q���?����}���u�f����\{�z�F�&��kT�h6!t��*|Ŗ�6�ݎ6�Ϩ����==�\�H����w�@/`�6}k����q�|p�����Pi{7Ba�1�=����ЛE���D2>�S�y\��ZE� 0.KgS��v����W>W!���55������g8���D��%0th�vq�b�6�� ����� ]nj���%6��)-F�g9w�WG��T�Ջ{��l ���0�\VSc#׷�eΰ"C��`h��J���P7�U�@��C���M  �FB¤�f�ewk/�;��f�\����Z�a����������!.�z1A����mFV�BB���T�Y�kX�� �{�TYc���0f��qv �Ri�{���>�8A�*b�]�S��7�=�~o+��c�7;�����'Y⩴��@�}~8����L���g 4�h7�g�+��߮���i��Q��CyWYq�e|�w���-By.�r�xB���<Nf�MV��?�����SK��ǹ	E���M�f�q�HI9-�U�2���Qgǻ#6��j�uo�_ѴAo��/�O�>>�n�	�k�Z��D �!�Ǎ��ע4�gc��E��Ņ�y���5[&���j��^-��f&���3/�VQL��$����P!�Ѣs�S��)���P3��_'N_�!aSl���]���>ey�7�\�鯋t����ʒ^��
� ����a
����(��lT����*|�4gD�o=�+C	%ɳuA!��IL���Ō�P��m�<�p���V��'/��ܳ �a��S������X)�81��n�{pw���^��e�{H�*��	0�g�{;��?�
&*��uHƊI����PCuO�7,A�{6%N�ʜ���(�����?Dv�	]�#��������d�s��h��Y�aivaM�0ɯ����]�d9b_Q�P�MSU��jLl5戥��h�Ly�۞�9�I�t����N���3�[�	h[�=��e����$&��O{���r@J�ɷ�N��2է�U���<�Ƒ��-����A�Q��L���I���kW�{Fh]���L�-�-���B}e/"���X�{�.�Q�ϊ�E���<�&�HU0y��LY@��rl����mQ��Fgz�`���5��H����6K7wg�KX*��*�=���%3�?���y�C_7��.�m�b�I߯a��v���q6���R#��J��$�`�� [��[����a@�3��X��e��?/;SG7�{~u!��sj~^��Q�Z��U̺��$���'���W�4ƶ� ���r�#D%�35�ٱ����f����	R�n�G��u��=�⒊w�"~��e��0*HX����#H��;$���W��܇�H`��Z#Q'7��`��Ъ��T-�I{�y�J��EO�[ec�pRKg ����F�S�F&qLlfJ���z�W��V5��Ebw}c=7vY(܆�8��Sz�RU^n���9�a҂�
�4�M�`R$)O�
/��p���16��0j �KfP#b�ML��J:��#����C/h��1{�>�Vp+)�ɏ_:�/8�5�=tw��i�4�O����y��+U�y!/�_ӣ��򣊂�P���Z��ynԻ$w9�~��U�|�V��'�
>����%��XR�����@��uA������r���mTC�-4�uec젍#�BF��F��2���.��C2�X�������7�o]�̠9���wt+�=��
����%�������f��-/��4���fw�{b�ag��cD���n�����M{���cT�sv�� ��)JH­i�k�+��� x@��D�I��j*Y��i-�[��,:��[�>�&��͉l��8@���Nh��H����8�˴Gt�-�
�P�g����\�\���s8N�[�����!�i 1��! /���?h�J��(5%���4%:q�ųvX�AE^�����2� �nƴ��n�lOEq<����N�f?Ӆ2\)IV�g���{'�y��"MD���iNAa�'U�}�=�����)�}�5�q>w����|�\�!O�1yG�Y<���L�	�8�Lk�׸�<�w΋n��͛P��Ҥ6�Y¯[HB<}��3����VOR�F9�M���i�}`���
3g�*���z/u�Y�nC����!n[�	}���B�@��^8�^����}p�:U�~� �gok�i}��n�{=����f�V�R)�x�>���|:++r'��^ŽIB:���E:�4�<��!����~u���i ��GY��J<��9�i�=j�m.��$#±��5�
�-S�o/����#�bd	������v�a�o����r���/ȇ=�:�r.�5�5��{�U[x����$2�6��#@\S�=e+��S����4������9����Vw�j�0����?�C����k�PA�*�i�q�35�������s(��A�HrT�/��ͪ��|�}:�y(�Zską�Y�dh6�<��:�ю]r*�Yօ��7�Q�2aBd ���J�FF��:�,�(��i����r�MlUO�`�b���B�Ls�V�~M����ި4�0�M���2Y%HR�m-��˺:th�����ۢ�q}.3����8b˗h*����%����C�C~��3��6ܥO���jB�=d��?7��⼹'�ΫS�|{���u��V��	��BF#�ob�UM���N�Rr����C��>�@��3�j8O_�F�Œ1�m�ޅF<жM�̡����Z��[��Kk�:��ds�v��i��NP����)��<#6HxۊY��QDk��f/�[�R�������²�9� �Д(~�^W��v7Ҕ%R@r����D~�D��lc���6�*��M%Q�`�kxx�[?� �ė	=@�/�3��=1�,��4��mS�㎩�a�A-��si?Qs`����߈���$x
'$�>�v�-/��s6��&EPZC������)��8D����(�/5^CԍD�#h�6�qB3�E
�7I�KQ��{�G�A7I��5�+}2xK$1��J�N)�Z�Y�X�}�C���Qoa�LQ�E���K��_8~��RTa\����+2��!*�ۼm�6�	��5����Ą, #�c]�I�vr��eX�3�V۴�8T���40�̀U��)�A��ә�遍�h�U�=s[�b��3����w�U	<&�ܖ�NV��A9��@+Z��څm˲qX� �Mfp�>}��i*v�C��T��wь�շ�4�q�}�g�rt�Ê���m�W�Eꡗ���a�Jz%�>	1F���xn��F�L_w<^!���e���V%|E�ugi�|��}{��Pc,3Bn�S��d�I�U�����o���m���D��d�&�N͗
L`�1���u����z�GCo�U�_�3x��O(ؓ�e��,;��77�[DՔ�Y�T���W�����j3W�U�������c8{؜���GN<^�z���d��rd��^�*�v�����ba�%Ӥ N���0l�Jc��"��E�P�D%P���e�51͹�^;1��i��[1������0$�p��U�9�-;?^bƧ ��ȥw`y+LC�� ِ���>i���ԮpA
s$)�4��V�-i[.ϫ� '��Ԡ�co�ΐ���R�UB�Q��~odI
��@)I�L�$;Z��r���\V�_��A&x�<H/%G���`�+l��X{�u�;H�1WQ�;�7��<��ך@����FK���6��t�9`��̵PY�K�n?޹i��r��-$����("�[?����B$y���o��K��)dS�K����ۑ-+��:�B�`@��x�;{��P]��(?E��Q,�A�vN$��~@�%W�a���wUT�.ۦ0;EK�,���H��l4����AȚ@�˘2H�̼����y��)!g�Iӡ���\������i77e���>|f6�d#MY��ЦM�&�Ny��Ǵ|�o���!��u�2�`�����Å�S�s�u�����W������D��-g�{����&�c*�.��L%#�tʥ�s�$N3PJU������#bV�P]4\0ڨ�S���Ke@.��7F�����3d�q��������B�3y�w:�¸�	��;��%k^����DD�7D1:��������ec�o� ��.Ş������GZ�O48ڒx���-���p�&ū;��Iɜ��s�	#�����b���P���J��xbG�N�O]���Kn3�J�uR��\����2cFiΔ��c�ý�a��pV!�9�Ӈff��nY�)M���y�W�\�4
� ��E�⧘K1+��+B���ż������P\�ħ[a���ïv���	��N�Ovd��Ni�Һ��T�s���z�����(�ba\q���uk5y�ƃ��`����Va��y4�������r>"$=���iB|�5�/����c:�`Q���qW�#�<"cm���� �������U��	�+G���qܘ��;� � �K��鵚ŭ��c�s�*��ۄ���S��*�O�d�p+Gu�UO'x��$*����M#��	�A.��a�1�kk��2�9F��T�����]a�K\�ZL�a�+�!���l;-��ΐ��(��@(�.�uN�
�zz�s�"ڿ�a����aԅ�Ej�g�P�!n��1F3�7���� <x�ֳN�ySROόbF@��.\w�wo�ʊ�����F����d�&�h��(��6�)>g��,�n�B�͹�}���=�5�������c_�����w;ꚾ��aX������A�p���eLs|�ڨ� ���;���,�!'�����B�~�w�W=�N
Y�h��	'��̀�,07uo��lW_�v	1��&�-�4?ws�����Ƹc�|>(7<Ж�$e��!��5�N�ms���>,@,]�0�A~v�l�]�+>^kÉ�p�D�j귎sl��u�f���@a��x�vQ�ݮ��%V�J�35k�2׉
�H�,��-�FrZ�7�U�q5���s��KbםdȞW�t�+��JX(�����K��ط#��{Ӧ�;��Ѭ�U
Se(�����_]�{$��������1 �}�w��k�}�v|Xb�Q�����!m��_��n�?�@�8u�i1�F5́��#/\��P��]#�0_�$��4�m�y�.��H���!��ؠ^D�ʭq����=(��տ�Oc��6�%Իh�@s˗`�YwY���0bg�:�-��$m#��5��_��܊���U��!q�>t�$&
��tZ&��ޝ�O�D�//�:���i[%ޮ1j�p�X�u��827؂�(_�(�ҚI~�F1K0x������c�Ѵ�3�
t���V��\�K�<�xӚ�K-�;m&֩���a�X��3k)�,4tm"QR{P�L�ΧlZ�ǀ��������"UKՅ�N��U�����CA���9$,�������nZ6�^m��[
��.�o�
���C=�'��E��4�m�m��PZT�T�C�-�>_QM�Э����1Buh���al3��*ot�F"A6AME5j�L%S�-�M�Y�4�pѪ'���C�颕�U:[�=@��ӄ#�o��rr�?�n�(����f�5�f�t��J�'��C�ޓQ���I�vc�,ٻ�tԇ6ӟ�&U� c��j���M�`<�c�{����4)#T��a3��
r�b���+"�ɯ�ޗ�w�>F��T����(���wf��*�-q�N`Ȼ�Le��ڠ���{'%����`�}��:v\�1�F�5���P�C�E*���;��z��D�����D���s?65?���/��J'Xx;�,x���O
u(gAj��s��኎@��ژU�Z{��?|}N�X�/\U��J (y�Q��@ù8�p���ћ��ݍ6�nr����.L۸�~�rb3�A���w��|
���y0�/Z�B$�O*
jKD&8��$P�<�l#��צk"�vJ��H�q2�URZR�]��(�R��N�I�W��d$�P�<X�<�Ľ)19y*Б��;;���?xwHw蔉�?�ӫ����?��z�d9I��dQ�����:ag�����:}���	_j@�3���|"���?�L��r����m������C�,�*�i�;��Ŝ�;Bro�;�*�<ӓh�lrۇ�_z��7��$e�fG����Z��KT�_W�^L�����X�v�b�?�t��L��������/��ݛ �^6ғ��UtE�cnX=��s�u�a�%�v�M����ð�p�Vd3G������<�Y�;���S&��A��wƹ	�@��9�!�R�T��8��=�K��p�:�g]��t�Ǽ������0!��j��g��rmkט,����p��Ls4�`�ҿ�����1�~�y�LS6������=փ.��4�g�D9�ő�e��Iqq�����&�1K��]sa*+�$�E�c2z��qߪ��P��_Y�e��n�%"t-+��ׯ����:��7cB�()Pof��_q6jV��>�Ox�3y4�Ne��}(?J���=��U\v�Z5�c����_�닻ֈ���o
����$+���' �����_��D_��)��f��ō��,c�/=>��qD-˸}HC̛�\��oz��F�b]\�9��W�ǉ+:�ܟo�!��/�o8���'�f�NqA1�Xu�m�����yf�kjR>.N�4��_��X�s�V�C2�>�{�m3'(��"�)Agh ��۬'X̘���N�¯��6��J�`���û;�b5������?I�[A�Lkq<�3\��X�ߘT[����F�����̥"Y�,A���g�&��C�e{HK;ۤ�2)O�0S��ᵒz�7��Lβ��L��/�v*���r�����^��명mo�nlR���!��)��ǉ��\P�\J߫S���T�ȑ�	��Y|���o�1���L�67�Şh�>Lѷi;
����~V6�f�j���s��n �Lj�OSU0~�����2s����JT�C�*МJyl K
��-�}IX��$�O1��x�w���҇y1�.x_�R@#J�n�3�<��(�	m(		bY}~P�Y7�Ό��!�0�ܽ:Å�����˨�^ns��M,Q�����D�����b�P�8��`�����&��O՚�b��a�:(�{Sh:��+���������}�$^��Vyޟ��ޫ�������cU�^�.�/#i7%H�T��.V�v�t�J2�4@�*l=]�\�v���1��� ��z�h���DgX`��u��dx��|��9��b�$��\�h*����B�#�̀��A���*.��[t��$����jez`���Wpc�G�Tb��S��������sw�Z��d_}���k^�2^����8Ј�?i�l�B;W�+q0O�Ql���M���y�/ơ毜K��Q&���y�v��0�@��j$#�{c���hl��$���@�=wF6��;c%���?4Qab\ӻ�����v�m/\���A��M��knJ0�óA{�s^6-�d���v'|�Ki��t��1�G]��JFKYs�<E�':=�c���3䲈��@!hB`��u��̼q��5/6��o���������6M�}�w�PJ&�Ό����(kmmᇶ	�	#|KAO����=�	3>������i�����	����rQ�P��u̺7�����3@�P���Q�o/SZ���`Z��M}��:�;~ޞ�����
����o�p�Q���hǢo���l���t�at[}��+�|w�8�p!A+sp��Pag[:m_0"�eTL(�Z�o��i玈����Ǵ�r��-�U2�T�����x(�g^�w��1�y���Yt^�{G\�W{l�%0<���T�j��[@f�Sɯ���P���x!g�����#86m�%N'|H���dH���#'�<yxx^��C3�,�k������G���Ƶ���F\Q�t�FFq�^��#0�1fV�������m��?b	�z��ˡT+ntX`���ț-�Sa[��ŹC���q6�[]|QnoO	k�\��k��y+�����`[�`N�m�z��d(�\�>�F���(���hN��P�[#MV��!dallx����%ȯMAE���8]�>��I���R`�>ߧg��	�]\�)�h��!;����\@��|���XfK��/���l`���m�@��50| 栎<6��­���̰�]��]���C�z#>� ����Rlr��A���%�3��XuA�����H�
/atZ�0v���P����	1�ݫ�ֳ��P�� � ��{�Mz �>�,9����ɢLX_��x#�N�/�F+Ff�(�}�b�)��8��-���-[Ջ��[�"�	��9  ��Ŋyvlp1g�U�	���l@��E�Ƣ��.t.�GX�ռE���|3���v�FIRf������#Իm�(��/���\�ͫn���d��/A�3��i,�Ar1�+A�X�H�86?"l��#�H���ji�_�6|���>=�����Z���u� �-�cۣG���$�~@����X5"c	�S��>7��o����C4�/LO�s�����[ac� SV/�qP-)��I����&�VG���(��,�����H�?�<
;�Hڧ zRȆ��YJ=b<w&�*�B�SB��x|D<�6 +p�G>��Ӌ/̶C�ZP~G�v�0����zKk��(s���R7�B-�f�{6��y�v�%!2V�4�f��O~��h�(>�V�~�*a?����{�zG��Tf�r�r>�*�Fn���;�t����T��r�L �Y>)*DZ��a��':��(���1/|��>G,P��Ui�7��XY�[��&�1-RKYM/x[ڥ��Y��)2J��ڛ6|���nhS��h��h�5O:���3���JV[ƣn��#%��\�^T�5T`,��1��m7�g�Ig�w���q�*��zPCu����&c�\A�*3G6@�xϡ������~��u��D�SQ!�+UMqKg�]$;Ztf�6�����T]�.+!w""2�`��q�}����?k
�h�HX|Y/���μ��_-�г.�5����$����K[i��:L�R��J���Z#�+[�9���[��ֻ^0�	^5���&�<�v/���H���EXv=uJ]�� �[���6+.=A�����7�Ȋ_��E	�XB��G���公�!Ӣ��]5w����!����N�����~�P&٬���Q�8�a��y���@k��h.�ױy�n͙.0g��L��S��0M�$��ի:�곦eUF_�m�)�j����ݟķ�#�b�{�Å��M��qc��w��6ka_�m��)*�?��_����1�e�I��a�͊�2��9���b�z�p���zÛ�9�$�f3J�59�{X�=��ˍa�{8�L�E��]W���(2D����#��(��{N1�⛏e�Oь�I��� )��v����I��:�CRQ��fR���B红�K��#$�	Z��p�V?���v�ug&h��fc������2V��ț��v��c\"s�I;vW�͊Dmq�u
.V�?�f�����4�еX��b�Hx�6eƣ%��:��L"�;�S'��\���M�f��w�S�������8DP�Bx�l�B�^��.�.6OUj�fO���h��&�&I�BF��Tc�L��I�\�1�j��:*p��G�gT!�qQ�D��ת��2��p�5\9'�e�w�X�E]�����#�2���,'�WT�6��đ�q����zPӳ����뙫��#�g,�^qy��_���8��������1�fvu� F�Мy�����r�ߞ�I+a�'۸���"b�^���^��.�T,��[����!j�c�q����T�Hb�H�9�.rl�6c^4���N�w�XgS3��ШR� �/��#��Iv���o&6��E�k`�}��h���a3ԗ�]*�L�ԁ�c'��R%NV���FKŶ��ឲ���Bh㺕���}��1VU:� �b������J�;xp�V���~����')��5�ɼ�`�X�q��R,po݉���X��8zBM`\[��!$��I��?�bM8b�Owݚ{#�W�\=z�n�(��XV�}��כq�-穥�M���gC�.C�M�r0!��F�';�>���1�L�]�;U0������S:��O=/�*�'1�%����[�G-��j�m��{v���)h�WĤ��8P��g�bk�3��v!M{�Aa@i���ٝ�#���������&���/��ۨ?/^P=Gma#E����ֽ_ �x���]�tR���U2��8�VB��i\���V�ԩT�\�`�gc�ݡ2��RV%�-j-�!8��Nِ��A���r���V|�!
"܇q��բ,<s#.�6�n��j��@��!�����Z�s��L�*z�eI�]υ���0��p������YXF\���Wik�z���
%��5��I��Y�� ���6�0�{XC'��0`�'@�^�)�u٫�7�g���-I�o߼�,T¾��.���M�k���*���E�c���1Dg�P�i������\9����k[뫥��'�=+
5�[�$4�^�.\־��W4��b2���o`�J��"��f�i*kD!�?*$ZE��v�m��1ȋ�S}oYDH�T��+v?İ�] ��J����~E�V�N�n��uS�9����jvqZՂ��)�dX�^ wǍ��t9c��cx~u�1X�b�(֜I@��otwc���G�P%e��и��T%
P5`a��E��c@)&���7�zY<V#��g�O��𬺺��-����>.]<�r����nͪ�p�.��S���HZi��v��j���Kܵ�f+�q�f����J��T���}V���ߡˡ�/���42`5\a�A�3���d�'8l���g�'2J��d����.�&t�Y4q�]�_������2�.#���ǖ�����]U�r�H��U��<�Հu��no���rJ�I���V`���?���{m��������{!	ƩCy]FE��1⢺����j6��F�=c�N*N㇘Ɯ\!�����^
��U� �W��[G�i��k�|�����������%/UL����lu����?9���Q�Uza�*
�v�Y���j�x��� �<+�.��>�X:�=GW�3�=X���9��A���b�Uc��;�19b���x��BAR9�H �t
i��&�0�7����X}.�����N����dzÓ`ne���2{u<���JdŸ��Qi�ps���.�#l�~>�k�Q[:��,N�&jw�xK��ě���^�E�8���q��+y�K��]���O`9�C�>�-J�S7��=���<}k�"X� _�	��@ʥ�s��
a�/b���)g�U�	��^�߀���;X7���6G��C̚��<��ף���h����U�.�{��Cc�_��!���X����?LsJ���NlE�j�K�-7$�>8�����~���p�^ê�	d����%����g�c>����Ge7��WxQ�n��I}>uBT/��,�x'���Ǔ��p<���fOq�g	i͸?J�
|�":צ�N���,g��1hxm��:��䢫���[���� aS���)�R�u\/��IbE�*MzJrxe�D��l�z!u*�ի��($�+2�]4]Quݔ-HM�/؂-��\Hy�=��?p!pu���e9퐔�u��)W��׫雯e7����7�H�w�{[��Ɗ���Ʉ�Or�����Ղ*0YBN�p�y��% K���v��C���;|��XQ���F���O]�{Bo�It�+��ڹa
0�mu' �n���|�
kEs�_��Lq2��̟��1�8nT�����2�L�
������	(�Ksv��S�<���!�PiS�t
�E�Q͟�ڶ�y^�.�}���*&&�j��Er�ݖ[ĶȔE��@�C9�0����Mq If@��%�fc�u��A���r���K
�f<@#��zAgJ��o+�옮�)�pq�����`?������'A�z�,S��2HFX�~ ��lŽ�L�m�%DX�[�N����m[S��>J��Ξ5����@��ؤڿ����aǛS�G%��ÿ����|X���O�S�
U-.���n�K�	�q۪�\��ښ%4V��M�-���k�N���c�!�Ò��L�z1���g?����q�sT�l�a��11A9���ށb��9���?
�:�q]�4e�,�hh?5��!�����m`��\'��F{����R�k8��B�FT��}��f�/�
ҷ��f�js;#���~�e������f{��zm�/�&���,Wv�{�k<a�<���;�Mҍ�o���g�<�+	��7�]��NM��k}�a\�J�����y��v}��``B�ű�3����}���m9%;ëP��P�o���/�{����r�1�M�P�O��G��YR�-�{KTUհ
޽4��!�Jؽ������*��6QxM����F�g��`�R�Rݯ
���S�c�Ӳx��>���Z��T�ܙl ��3����}�pe�\޶�+�U�HΠ��ErQ�kO�+a�*�����"�tm�=�SBd�I&�n�
�`����cԚ����J�i��]۾�%J�i�D4�z`�hm���D3�Ť���>i�~!�y� �Fn�b9�i�+�q-��@t������1�[#��z:#!��g%4-�*�X�׾�E>�n#=o��bfƟ�z^�N՟�"�dkO@b���W�F���]�;OA�q�2V��;�=��,�Ԗ�Ձ$J'Q�U��-�>�!A-V�
=l�x�ܧh������Tj�F9�9P_���2�%�js�f�۸��3��fˍ�8a�v*l7-߃�-��L\U꺏�^!� �z�ZuT\U] �\e�UD��L���1WH�V��fm�w�� ���I�8q��F(X��� ���_��*b:�����vR�Vǁ�/�X)�S�#��c���PB� ����{Ī~�؏��7�����4󡯀�p���S2�QV(Q�W�\��ׯ>��;w�q^�]�~�K7���F-[3,x�~"BI��͠�%��������Vy��6>ѦYL�6~0D�~@�7ƧBp��:K>�`��x������rE�lF�BNs�?�_X�w�s����!���{7*su��mU����.�J��Mp��e2N�p.Q�KX�חQ��!4�O�(,�����b����)O5��_e����^'Y<K��������Z��Csy�~�II͒DlS{�`̳_��!�8j���BS���Xn�Нw���:�3a][�r^�0N Md��y�G��pm�� ���#���i\���Z8����u�P�ז�Ž� jF
�ŘN����@�e�/c�T�}*��|5� w+�X4nIp>��J}�G�o���;�J**���"��c\����Xߘ�N�݇p;в�1����O%%=u�0.��z�z�_�� �wJ��c�]��V~�R��!���8_�?���%�b=�`h�{�-����t�������[[<0�h#�2���P����yg>M�?��Z����k� ��N���O���u� ���Ľ��x�*(�\��=��t����ڊ�**�-��-�mL��}1�)}��y�I�}�^U(VFd�8>�56Mk���Ʃ*?+��ݍ�����+a�ŷ�Ƈ{��w�����g�/���j�$+8l��^��:��q� C�|�(_�N{���K4�����[���9�0��ke7E��UB�(7����4T�h��x� �M3᭦D��N��>�GK��(s �/�+ﲣ�����.��E�j�$���u'+4��O�u����P�	�v�v������9�"Z&a"�SU���K,-z��W�$�^��*�qj-��+77��x��T�gֆ����9�5��g9��zw)��� \ƨ�fw�q��7QhD���PKm��h0j����৤��u����\�XW]E����8 ����̢�(���A?��>O8K�N��<ֽ��¶j!Z��Pb��x��Y�?�4��Gl`�ٍ�Y�BW���֤Fm���o^���4Ψ ����->ؔK��	x��Q#�x4�#p���9�����h�E ڶ�p�8�AOk=�H:=>�)��f�MI\�C�D!!�|mUպI y/��x��BA[�� ��3�[
f�٨6�U�&ǯ�2[Z�_�x���~��<yQ!��tW���i�?�5���!A�'��!D-�­������J�N5�#��}�6.rS9���=���^���(��-����{�>�]�t�M��ʋT:J�	��|���]��b�8h]/�c�S�Z�K���W���%˲s�'�g��8����*���d�ы�r�8��ln���A��\H��艎�%�N��I,�s)E��w���_I��uR ô#��h�]���
ެ�-��X�����h7��S��}	kx8�d��{����c��K�����;��������v���n���NunF���E���� ���3�ws�YG�|LNאD��5�y�n��=�5u;�"y �w"_{��<��^y	�C`���+�$��	-�,�f�����\󞾒�;����%޼dL��M�V}�N��P'�4���w:?y�C
�a<�� ��?�w3���{��z�.zjc�.!<Q����T����ի��,L^W�%��|���a,H�]ʭ�G
F~��K�L��n�)��Tk�Jr�#�WJ����Q�2�M��0��e��h��	_��}� ��[l>��̗�a��
S������ڀ���6.��hzr�.�tؓ�#ٴ�5,L�k!��J�ߗI>�-���%3��?��C����1����"���I�7/�CI�I�wU���;Z-M�����~$�%��1��*�m�T�/�Dv��N	��s������?Ǳ~�o^���fŏ�[(�Zfܧz�����=i����}��q=���'S�]�=��c~6r�ȉBb�f��Y!�*�F�Snq�3k ��r���O��d��M����_���ՂA����=h��8��q^��Mwu���f2���ڕl�ZȰf�~�{���� ���9L�-4�iu�Rn[�ƺҁ�Z3�'�fM�&<�t�-A�*���pW��L�Ӵ�/�}Biϔ%0���8#Rlg|�P:+��xH�~�a�Ͻ8��(��"B/#c�}���s�)nr�E>02v��L�B��f��U�o���7a����rs�iS���@���~��Y���-����8���ۊl�}�6�,�՗SYhƷЖ�n�3�%	^����#İ}lu�?����-���xk�:x�^C+�H�,{ў2e��tԍ2Npw�s�Z3��(I���m
%s���+��Q�#��@zl�_��MJN���pE�&��Q~\X��Ko�FS35�����M-p�����s7k��?�;GFP+����9�OjO�v��3��
��4��1	�t�!n1���喺���J_\����Rȁ��М�E
;r�V�=����	���R# !��|���L&sSߩ��_�����sZ}���g%<��9}&m��o#��mA! �&�tπ	�||����K6�>��4�W^��i���Phk�����ҥ�y1T��+����!_Ul�b]j�4����ö?M�L���{\ơ�x����he_e"���)��O�<k�(F���\��ۺ�}�$��p�`�*z�m�T��(D�aW�^�;q� !F� ˲o)ǃ��p��Hjf-f�9����j��q�^��^8c�_�)��q�������q089�#�#�cm��;R:�j�E��f��A�>'��ďo۔ .����M������(%!7G`VZ����4��]u�l_ؘ�vX�fk���-*��&vG���[��h��Q�Jw��1�2dƨNltU���lھ
l��4YZ������>H�������Wd�DU&��S.��U�ol?�:��x�����;"�я(�Ͼ��Z�[7�	W�5�%ߗsR�����@�K�F�~ƾ� ���-O�VG�m��� &��n�Zy��r�'�l0c��M�� DM��Y1���P�͎#y�*l�����@�`���~�VJjz^�P�K5�=��?�ޫB]�2�Q.Q�R�I{!�f8-�-n{5�=�������7�V�J�B��7k2kβt]�Iyk�g5ɝ�;_�g�
h�w���:�dUm���-�s�
J����oD�)ا��<b�晸�p~��v)��V��~��df����	�sWq�_�s���<-Rm!Zu�bQI��T�0|3U��Q���T?�ڟ���=��"��-�A��N�Γ�,��B߈�s�����-|�K�>%���+�9CTc�S@�t�@Z+�`�{M�/&d��Z8��83�n�r=�s2�;'� .(����x��e�YY��FD�b���i�O�fB[�j��=@�v._�� 5�k�:�͘����Y$��m���U�}��=h+%fk����C_�Ȫ��pI�Vf,�!+��΍9^�y������aB��hr�;驜�Z1^ɹ�~]�{6���Ӂb�[��a@ �ґh�m+%�鷞r�_-��$����i���}D�،�H�ʊ�K�eň`͝� :���fl�aX-)�"PZ�v8Q�+���Hp�:���"����
��s������x�f���#��=�	K��SϺ�Һ��\~d�M*Y�
�	k�񼌸�NT�>`u̐0o��Z��J{�8S[��oK�ٯ�Gޮ�\&�`���J�G�u_a�?�2d���#�>�l4,�+h�h$u���i�N�x�ԩ���{�_;"Ӱr�EܵH���gdn�`�����JUX�f�C�k��$i��k�*��İ߱w���j;�g�u�tw�K�YcV13�g�̝�C%7�5��B2vg��
�o�ַ�/~�&u�����M{(��aZ��*��s�zK�֛�U��p9�T��o�����Y:\&�|KMɉ�,Tgk5uc�����5��5�.h�R?n��h$�S<�O��i�� @7!����$���M?e�E����}A��4tJ} w	�>��WW������f�Nş���(�H��r���a�B���%���?%�]�I���c�4Ak��/S�Nq�`vS�	�%l!/�lm2����(��B�6;�bj��J����^���[v}dn�d��d�4���p���O�zu��+鸡�6)hf/�Iǌ\z8B��=��R�4Ҥ�L;�I�d��Ex"�r֨���_��
��F3n!�������|}�k��ei��q\���Ծ�R��&��UO��w���|j��SG��x_ 4�e���d�i<=Z2����" Hk�J�0��c"k�F p�0�Y�B���5��P���XX�٠Ĉ0e��	#뭳�2T�}�lvS�'�QS��R��5$nޯ�M�bu��C�+��]�\���ϟd�g(?)c)��*��9�S�z��.À�N�7�nJ�L���卜���5h�@���ڵ����.�~$v�U�XS��?v* ��k�ҫo�d$Ʈ����V]Hn/�D�*Ke��iWb�gUs����=��o�u��9�D��A������'�½/�.�	����M��*���{���vdӌ$s]\X3���Bk��Jm?Ǻ}�'?n'(�g�$�=C�\uE��Z0&�2R�]�C�ġ�s��Sb�_�J���E�O�db�Hk�
ξX�i�˙�:�;��_�J�.A �r�r�m������pJ����/�A��nZ��b�b/{�.<K�U.C,������,6~�!�Z�V���u�����y�x8�\�ҏ`���S��<s�b6��<P��o�pcq�|Nى�AmZ�7��n�ik���D:��{�ϳ�b�������ǻ�c�B;ĬXn\�!����"�~�V��t� 6���/n�3����m>�r$b�t�,�M�x�.����]=�Պ�|̀��zha"ї��KU�e|n��T�HR]�Q��:ҵ{ŋ��]���A=��8��^��>��E�tx�K�Q?�B/0��B���J9b�3_�J����ZӲp�z1X{��e�i:&�)A�o� Y-}R���npw�JJ�Bdo�,��øՆ�(t�.��+�~�8ٞ3^!�g� 7���9ڤqC����[X�\,��|���F��^�H~k	��>��[�3ҟe�/�P܆��*���\:N�5��o�?�>�uH�5'�w��,����x�}�@r͊g�߳�ⲷ#� �P�}�W.C�G�5�1�v��t[L^W��7����ҙ�.v������l�U*	�hy�=�.i��Y���;�b��@K{li&ѯ#Q��]6�L��p�a¿�T�����F0��G�#�D��bj��Regt�[�Q�u��;xG��a��U�q:��ov�LǘS�_��ijD�٬�1�jUE�Q��P��K�VbK@�dk��\���x�C*���0�����p���׉k��[m��[��G�d3�'��@��l�h��=�S�h*��p(Yπ����W��H��Ԕ\��#���	9�~��na��4�>���I�(�u/��J+��	��]0Co����v��������P��#��ا�A�?K�ƈ���c���#�] 
�pr�}��m����\E�!����#�G9۰b�a� ��V�o_�"׿zo����V��)�^k�LuH�E�Ē8o'w���8���4y9���n�2C�Q�5�o�{����@�*�A�ps�{s����2\P��G�b��r�<IZ֘�)�Ũ'�����P��ݤH��'��Q0�9HB���OZ��]�$�V�X��g���B�z��Pg��VI.T�ż�;٧[�rw��4���Dl�D�	V�*��z��n�?N�qX��pн�b���d��ʁ��(N	�\z�_��C6���o;�/�.�O�p]~�:InXf���;�ч���ʱQ��G��ӎtU�n|D����q�� �9�'0*Ҁ0�*�� ���j�mn�}���8��'y-]�^!�T��DRڟ�?��^��2��/�l;���Dp0J{>s5�-W�E�c"��8�0/p�}|b�g�s�<�����j�hT,M]���=�FGb�;�-����k�|o���'S$�t�M��_���:���ר�~�e�� �W��N����	Q����wCI2{�%�M#�";oV��K1ǀ���qgb�_�vr�e�,�7�S¹����R� M�@�6�d #�������B��k䁷���E���y��vZ�0+9r}��mYct�J"���سRr��˵��I~�n��(x.��3���d8K�2g�N�fBs�Y�M!�sY���xU�N�5}ҁ��?R�}s ��[��u;t�I���y�(�2��
��U�;,$	�Ӽ5�çLD	�*ĭ����d��-�V�ŢG�0�3v"��qc{~�T�^s�\�ֿg ��6��3�g��vS� -\ܣY?�m7/�m��
�ǫ�,C�j�h�;Y�l]�ńk��^4̃��S)��1����k�j�FG�U�@���u�׆���Ч$���Ć��T8����$�����.�Z �Ǐt�Ga4Uۂ�/4�g�.Ԅ��VF�b��$���*�K,q���Ca�r�G��UCǇI������߾Zz�Q7-r��Q��i>uԙ�Х�(1���	�ߣ�0ĸ(�cf5�^���l~g{�s0[�U	��r�/0���T�(W���y���Pʵ��>S�lȚ���M��c��/�0i��<j#��5���QX_8s!_5X�1�S��<�4���D*�����H�~�)Ad1 U�6�VU��Q��]K��]&l��$��'TV�\��/�CZC�.}u*��o��X��!�ڰ#�n#\���8�0;��: �E5�I��_��39�P���t ��`x5�눀���򖭒�����}������L� Z�{���jRK>�T���w�G��2��W�#L�DgK��s��r�u��(W}�aP�̳#4߫w�Rn@�C����o�,.��ܿ�֫�ʴWe�"%�}|�c�F��������U��x��d�{p#�v+�׮�c���0����H(�D]�՝�棗�}ߑ���d�� �XÄ�Wc�=��m:���3W����|�3�� >�gR�(��a���4���Ƴ�x}ٛ[�OJ���Oɡ���`< ��h4m�le�3^&V6TYџU����|�<��F�pP&���J@r���I��6�i�)w�|쟥�v~·DZ �}�Zf~����W�a!�b� iw� �h�����h��-��H���o�`��O�y`ʓ����{e
|�y�b�)y���Tk:�֢��n�zmx�"!�+w��j.�
���a7��!��j�����Ϭ��PM�p�xb�*4�lf���O�#\`�ʕ	�s��B7�<2�3��-��O[ŭ2A�s��-� ��cỼP����Ƥg#9.�O(H�ױ�~{]�ki���*P��I��j)*�"�m�&��*�U�佭B�p�1(�K���[DW$[��9±/�xr}�5����ZIP_����b�n�g��]Ո��*)gR���:,�9����;]�o���gQ�o7�j�k��y�Y7��Y�Z�]i�a��H��$� �4���暨7hʏ�^�`mɶ�)�I��En����;ۍ����.��m�z�J$�`?[<<o�ax�[#�������Óm��V�������@��d�QEKN�D�m1xa()2/�#����r���L��[� �
}���<�Zܴ�#Y�v )l�c���u���eJ��b��?6=�z'�မ�����C���J;�#������o^§K7��R�p%RG�[��Lȉ�ݽ�[#V�&�kI��&zc�����٠d���=�Vw�.ͼ�/���'�	�8!懅|�PT��.W���]�{F(��Ґ\a��y[��������ӟ!¤�gk1��W7��*aTI�>� -������K� �{���<1��w��|�阔j������\�}$������(A�܂��ޖCU�|�A�a4WZ�7y�BL8"�L�/��̓����Ee7��������,�@2٠�7�?��r9�H��-�_���yhݥ>�1?>��Bܺ��9|��PI�㎅d/����~�t���V#A~"�4\�%O�K��:fl3����K���i���:�FZ�͇�h
���.Ȏj�{��qX��$��úD�k��%����
�6'���z{o���0���������+��D�4H(�tt���@�)��m��Բ�J�t4�`�lI��r ?�P��sdʄ.H���I#2|�C �]R�D��,���z��
�s���4ti4)�#�F�X�*"v6�zL�?��_I3�/X�+	M㎫PM��3�t���/@���2]��P��[ǒ�Ȓʹ�X�.+�%g4<�H��%tJ���n�?�PE0�;+�����?�a{���̠���>l^����qt8�2v��@�!�.�Z�Ꞡ�T��b��ey�}���PD��t�ԟ��?�eTäG�)�llj%�T2��0-���,L�,�?�*�!|�]Q�5����tc�74�Ӑ�VBPJ���Y��g��n�2��Y����j�>����k[B'����d{�/�6�l'�Lxt��v=.�e�ָ���U�^� �L��o���U�gw��d�l3���fʽ���շ�#d�yY��Gb�5sD3$�_��o�����/B���h]�4��p�����U~t�h�6}k��\@^�7O	��1�����k&���j�� �8����2P�0bFfH����L8cP8�q�����Nr���#ȸ�4�X%��K�I]����L�N��r�� ���<�-�<�.� ��n�n�#�<��{K�W}\���N.�A����,��XRwok�2�,��6���:�?�Ax83��9G����R�>�io��I���0�ޏ���${Wl�p���x#�c�x�J�jT�Q}��ڈo	Tp��!鰐WWM��L��8!�d�֬���G���X�
i1����ꙋۄ���#�k�tW�B6�>�#W��J�x�?c����Q�%u��t�����F�/�jjN�%u��EP������B���n��xiz�H��~ܦy��P9�)n"�I����G�ɒ*j'�cS�\ߟ2�,y�1&�AI{Q@ B�%����`���l��&g���l
���IkTଚ�p%��4�5����W�Ol������Ste��1��^J�T�Ű���D��1�~�%��R��yKk�*�A�x �SZ��H�2�gtA��/�F|]�ɓE1�ne���}�ڜ��?GS|�[m���xԷ�ο�"���?8o�0�[K�	`�ޓk�3�M�6ݺ�-�o��Ep�����H/tK,8W� O\� �<�l�:��	����3�y�Z&bGO�E3ݡ���}���3V C�F}ȕ1�ydbf���W���?Ԓ��(k��*�
C+���L�\�=�����-���7B|]�/�#'K���<q�k��J7�O��{����e>Z��(:��V���<\/�����G���Ί�B:֜�)��}ߦ��I�|��^A��Bv��n r���b����![69��_�ׯ�Z����ԥ{�B���۰bg�$����/�1io�ɶ�F���-�>}����4�^��l+94�rb	��4������5}bb����E�B��fB��bv'�b���� �K���L��3� ��ۀ�Xc��t�ĉ�r�0��N�����Ȥ«
\��uB"��"
Q����P�������D�dvRW�ԶQ!S�wB;����{�GbN�^�G=������R5���c�"%��y�R4<��o�ǐ��(�l�m� �	:����|��p1O7q]���u;���w2�J͒��Ե�݃���`.���9x��Co��L���m��f�n�i?-�;��ze��p�h�n��CM�r:�sɭ�z�_�\���,\�y�qU1�
e��
R5A���)} K�Lg��&U�(<�@����Z�	�M���G\�oj�$#t�z�Y���y���	�f����=}Ku��_G�,���8	>om���2]���
��oo����i@�+\�+�I,r!ۍo*m�����;���E�K�_g���'2�l<����@��g�E5q�'�g/����I��n�;�����c_5=���o��qxY]�~�-��{���	�������[W�G@2�!䉿.�5�	��GY�2("�f)�.��Ϝv��trֳI�/��rk�H"��ɫ���܎�옎�S
�g:ۭ����p��E�b�$���>�:,h�6d\�֨����|����%T��YE"At��&�U�?�Y3���b��o1�&W��أy*�u�I%��0Z�����"<��"�.�D���y����A8����p
���.m��.xz}��N��[~�"H��PrB^�uYC���5�sL�SǶ�8j�+�H�Ia�� S�r������X���/<�|굥�� J4/D۶��G��vd�ÓB���D�v�
��8i����|������dr�gb � � ΀��#������ԫ��\,����}�������e��,^!s��_��ږ�WU��F�����|Cs��tWf���A7����}�"ћ�G{��1
�&R�W�RN�ii���|9��q�`��컠)�h����6�'DVEC�K�v3S1���n'�k�HV(N*㝁�sh����rկu�4�\J��f�>mbuOe�c����b �F2��I+?��E2`�&��C��k�)M8/�M!r�xk�iRG�SrK,pC����SֶA�$�<ʄN�^�u)`�@�8��b��2�+�x������چ��h��vr�P�J��mk�˟�p<4:��ʩj��W��GT���(g�ԑ���j�:૪��}���v��𺫺>k->�+q0ڲ��
h�ES�ټ���#�w( Ĺ-Mʴ�E0)�p�qf��������@u��쫊ZO�'�M����2�@��/���$�ɀ�`A�ڵ� i���Z{�{��Þ0��M��{"���f��s���mU3k*�g`3�H)B��
�+�S=���l|zj^���6������ؓ!����kp2�>m[��oi0���}g0)QJn�s�N�U�4������Y��������X�(~P͡���׉r.?��Ż�z>��� :ɂ�M\�F�S%��_T�ҋ��w������'�Sxb��*�T�Ca�>���9G�Jprќ�� ��a/ l�	������զ�L���֝�t�SG����(#K{�$>S���W4F9A����ז���A�ck4�g��+Ҷ_Z�$�>�$q!����HRDVf0%e��E	wȢ�.@1�}��� !�;x�I� �8�È������Ӯ�[�KP`XѲ8ӊ��3Lٱz�T�W��.(���;�˦2E:̸�$�\G�������;OuF��3���U"���n`m�YՕ��b]U�ga+ZĿ���	��`�i'R+;@@ޘ� e���<3�.��uX��tkM��r2x���ة�K��1�Q�h�mG��p��J��` �+-��'��7h`��Z��p�-n<˩���*2�՘������~�+��پ _D$d��b��̳�����������Fi��k�#jp�xs,�J���E��C�{��^o[��щf.?/�F����Y���K�N�`�@������A�,���Q��N��{q쌇%�����.,Z���q^X:ꈀ5S۴RU��.[���F�+�)�l�dG[Y�d����G�]}S�e���G ��vyB�f츞r<ۂŴ+���l�G�z;+6Wj>��(�ʅ��x�0�Y�Q>���q3�`�!{�v��I�񫂤3��<g�<�/��fg;�`$���I}�(PƁUL����A>0��0Q�]Y�4�����^.;�]
�xݘ�<���ϵ%l#G�(��u+��|Jξ=�K|��*�t>��"OO�x�^(���{.�r/���R��SC|��+Ʌ粝��6k�O��ym��` #�gv����ta�3���h�����[�f��J��͘��C��?��珚8��Y���vm��H��+jJޓ#.���
�^��׹a��u&,2�����X�X}�oJ1Y����-�����p~�r�:�P���t�Cb��[�dm8縃M�>��])>\<� 	�/b�1�e�	���.�S��Z� ��u�����h��@bm%F=�8�iIyƃt�"㫙��yt�×�:��V�'���
����_�p����`����������r���
�[Ì��`9j! �U��W	����fq/n'�w�}�*Z��"{�\e��na/�����	���
�Op���}��X�:��v3(�x3n�r���|�d�m�����P~z��P����&��l��Y��v�f�2D ��Q�J%��uP�K�9r_/�����V�����i`k�i`��NS�����\��<m�ND�X�g��?�����Ʀ��%h���cb�6905�U��L0H=��;;R���;\u�}$~5����� X�aJ�Q��P#����S��,�H�XAd�'E��]%�%�k����T��4K2��Q���"N�X��u�)����Eڵ�H�jo��jã��૓�}�[��Wl�\Z%~#E�<*�o1 5$�=D�q�n��¸��jX��� w����Ɉ�V�����d���L}��5YF�Yg���9��Z�A�H�!�Czخ���3n%����b�Z-y�*a� A��\BſLP E{W/�����+����2*���_0Ƌr�W����N�BӋ;��e�qrNP�NqaOC����@��~�C�����`�Cm�����PB�
&>?ۇ�`��C}tӱ�իz�΅v�F��T�Ӆ��Uk��p��CA!7c{`oʆ�>���Z���䓈��X����~���E�����d�#1}�4n�ⴝ j,��A������@h����d����M_�C1�_���J.2��/�TJ��M��a����?�FX_U÷Ӫ��Yd��W�~�L5���A� �S.y�X#�wh��O䖵}||�/�`˳'�x�14	|!����ꄘ�E�[ϙh��ڮ)#�o+��@�si��1�j��A5�E��O���;�-�F�YRL�>����x��C�VJ�Q�I��?���%(��� �����U y.�[��}��l��(t�#�B�,��� �u�H𮋫&���g@����40�mң�M��l]ك-zy�ӄ^�~��K/\��GE�D���L�}�L��q���K�:���`�-
f��U��@��?;If��3Jx��`��̺���Q���Y-��_okN�\�H���B-m�8*!q�t?�ˀ������������F�HL�A��6���,��K��w��fLA@f&f���H�u�g���_�=�^`�Ir�o�ux+R��P+�����K[���}),'�t%�y4,R�BI,y֡.�[���Չ���B����Jp�?D����6����H��� �	[U�A���{�F�:�TگD?)#
�I&o��u�{t	g%�藙}�fkᣥ�E�.��QQ��9�΍��G!u�zG��;[5��	h0.��-�wr��m��i%^�a�4 [8�r�6��n3SH�޶����ғ�z�J����ϐ�؏a6�o���v|m�B�;D$U6�2��T����h3��}�p����t�~q}"����C4�\�U�PoZ�a������(�3�O��Ը�V�7qan;TK����^
n��!���&M ���T�VV��E�^C0�A�����D�șMZ4��EA��}B��T���Q�1-�8dS��^ga /���!>���[ɇ����ʴ$�13���/
a��<$Z�e�";��|k{!Jm�N�Y����8�0��ZI�C-S�6I��``��E>8��`�1n־���k�H%f_,�T��5L�VXh[��BQo��|�FD{�VM��}�3m�$w��{� ���s���µ���Ţ^�lDo�g�W��QW~��k���KX�@�����#����N���Q9�]r+I����5$f��Bͷ��}�N��7���Pu#�`��~�t�����n��Kh�q��Bw�$m������J��in!���W��z�S�>�:W�$*�~ `u�O��k�yH$�w~���+�����PHU[�ϯE4�gkE��?�O@�j=����.�w#PO/sy��o�y�#^U��-G��f�j�Y�ww5H��O����sQ�;M����|�����u�=oo33�<0G���ָ�A����g,E��y��uqi�����O&����(	��Lq�z�/��T�f=��6����L%U�A��[���	���/@uL,]�?^���?���=�q��m��P�}%M�P����Oe����O�lv�{�os���p�$f��/���`������my�)�埧�U$��1|b/�������	�B1�;�0��,�5i��������N-� K�q���4븻���t��?9��R��H�+�
l��r��!-�ar&�m�v�K=��͔7���/˂������<�@m��pA�T�,Cٽ�4�2�����7�e<�F�` �ǏrO��$��n ���#8����KAc���C7�.+M�߯L?�*�wHl�)��}�$��v��-Z6���
ҳ_�G�I��a?MgYG˓��e4��B��{������"�$=�z�L��xܸ[����U��Bp�PV��:�	�X\���Y:
�f�p�N�҆=���6�g�u�����A5��|(H�&d�_·�k�]��Nr4��I��n n1���+�����[��r��ӄ�b��1rQ�VQ�I�d%M.m�&Gl@�[�{�$+�B�ޖ2w� ����x�~y��5֏�y���e6m�\-S��~�U�!]ӆ1��P6~ ��jmGccMa���aܩ�U�h�o��!�\��1�΀�Q��k��rf���b4�L��J�s�&L�{�o�O���C���[�>;��W�w��d��XLwb)��:��T��>�0����X�(��F��8�C|��^�m`-Z��ynh2�P����~��h/���1
a�ͥ����B�mv�n+��+�SD]��
r�T�dY
�P�S�hf�ٌ��*򶘡��԰�:�YL|R���!�@Wpt%��,�ކL����C��j໑(HՄ�h��:��f��aCb��o#�7p_�}+J�Y��2�fg <w��{����¿�0�Z��1b�J�m	$��b���:n���_j�ͦ���2��0�D���#a�i�'�uA��]l���~ōP���+��9#�^���^;�O��3N��d�Ӭ9.���R�u����m�'������N}�W��Xh
Sk+Pqn9�r��t\�8�kz�5T��v�l����Z�EM��?�Mws�X6�e�������.�ԏ<8�OmHB�3��K���Yѱ*BI=Q����#V���&1��|�[t��F!�wҵ�)�anm	����k�W��z�u�� �!�/aA��7C��;z.�! 潊��wr���[Є��K�=��1�����h�y��a���+>!ǆsM9���4@��h��@�hPK�^T����Ʊ�Ev������|��0�E3/z)�5�#��u�Rku1e��&$��&�[�.砇̀|(;Ч;*'87��_��J�"��v@1_{�x����/����wԊ��[3����,��;�`�Ԩ�NB<Q���GO)���ʟ�*�)d���z��0��lUN��*�����Y�G2&�e��9�v��� V�Ag&�w�S/,5�-E��"0^zU֫�8R{"�T(��:_A��dd�'S��^�6s��ti�E,��H�L���r-f�e���	Qo�����z���:~#�&C�/����J�����U��Ʌ���xS��	�C��!(0NrՓ�E����|ZB�f`�xHe�S�R���r��H�+�8�{�aHh��&�E]w�,q�nB����R�E���ou�kz�#{V/>2_Z�.�5{�N�	3lי��f��K�e�N�G�L[�Ff���@x����
I�&�.Z�Amf�Th
y�������?c�Q���2yc�Csv%r���O���U٫H�b̋GΖL�����ft���Z���Ŵ�]U;��('`'1�6�8z���Aq����l��^�3��%��N���� �%��q{ə����y��\�����~Ҍ��*_P�&F(7�D"�e����C�N����jQ�`a`j:8���w[Si�5���xmn��ÖN{��(ĵ�Q�T=]P��J��?� [[��8�0�4���jP�i�);	rJ��QP$�����@y#&���m���I��`G����!�>���R����_�͓�����Vw�BAAa���e�����
�p�����ᶚ�/�	�O~����xm��D�#q�C`R��t'd�K�{i����ԨO�m�H��fa��Zc`q����p��f�f����md�*���3��9~0

I-p6�vVI�*���W#5L�(�4?�)�g6�A�A�ۨW��^�+c�an�=��?a���������yQ[�y�`c��Z��M{Y�"�� ;K�lŝ�@ҝ$�E�)�	����nO���#�<~��q�+�Z�1��_�M����Լqx,��4���|��J}��T[�����Z��'���;���Ĝ�̷d~�����m��`�$Xf���`����v���p@��M0S���bf���=7t���W�e�1���f?%D�F\k���8I�|�R.�2�=�xj��7a�j�߻6���):$r)������[�5�Ŏ����mjX/��ҟ�6ۦ�u;k� �e�C�蛂k�k��v`ч5PY�8f+-��fA�U����et0�S�-����f�&y�����[n$�`qɜM�4#X�(��|��!�a�'$�L�F"K�%�P��x���\�����p��{8�W���+9�-D!�b��j�� |���F>ʖ�;�cy	)U�	�����ٗ/�VVQ徫S���v��8\��I��M!��y2��ч�T�)N���EvRŦl��>�B�'�36ON�f�r�6�Q�3��Wez-v,�1@ЂBt����iB���t����z)�zߘ�i�M=Hp�7xǬU����F�X�3�d*~��y'������,c*��SD���QX�k�٦��h?��P��j_8�'�3-���i)��/�@1�ޓ�(03��,g2��+*w^Ğ!�Z�6AB������R
�Q6]�Uapƈ;�Q֦n�P(����;N�e���*�ĥ����d��W���1�N�g	�3	��k�Y�u�2�?�d�x�|��C�C��_b�钁�H����̑�%(���0ΉX��*4p��`�:i�	���;0��	}��_�~�R��:e>����^ͪ�Z�*-�F(w䶂J\�͚j�Π�[��ֱ�
Y(:]��Ѭ����d>O�s�}n�g}�����[�����,��D�t
R�����X��N���2S7h�n��~�\��ٞ,�#a{�D�$d-��U�L�Bok��n�30�p�!�2�����)�����"����A�8]�;��L�e�n�@/�>@�d�@�2qb��~��s��=Q/l�~��cPD��@V%f�:�#��R��yV�6�����X��0��Η8"��cn��L)�w5�Z�r ��j�g���>��u��)k������W��Yۘ����#��y�{��f��k�>��W�ۄ=:�<��aQp�l�W�~yE3�~�hu^��Z)��,�=zۀ�-�d��t=�d�5�-��N��g}��l���~Ab�D��$B[��Nk.k5ng�5�f�)<��,�oyHG����8�>G�t�P�mlYP�rˤ�5ج�������r�O[R�q���
?��u<�	(�.G�[q�dk'�m&�=Й�qZ)�N�M���4A���}I�{{�$��յn5�"�@N����1� �G!M��%\H)+���c��֯yY����i�IS��+%%^%�Z[b	 j��'3����O�Y�?k���