��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����gw���hK&,6�}x�Y�0zwզ�6K���<F^��jNB�(��ߕѦ|���+��3�UCR3�Lth�Y�ˎ��o]Z��y�����>���D�9�N���28Hd/��S�a3��@��!iW5�
�L�(���uG�����29��ruqV���eTX��""��v�Dr3V!��8���M+_ ��|�{)=쪩��:0���\8�c
�HD�6��ԕ�x���1o���~�_n�\�O3#���OZ(�z&	QBtA}�Ɯ>�M i���)��g��b�Y�?���ʹ�����r(Pz�>����1���Ħ��*u(�m�]sH�<<����T���V!�>��R@�
�_9���$G�'�a>�.��UP��~����.�?z�0����}��1�9����b5�����b�>��\F<�o���o����&���.��$%P�*ƣ͌YbVA`Q_��5f�?,��>|����9��Ǹ�S��}��RM6�+�3��Sp�+�FCo[8�r�W1˭	�x�.�%!2V�LԿ�۟�y
Nu�D�4ˊ
�b]�g��>��.��?�Nca��rs�Pڂ���-�ٝ_ّ���Pc�!iz:��,9G�L�H�.�3�o#�!�fK�{����j�:��Vﺦ�`�2�:����0:��������k[�!tv�Jn�i����y󩾜�v���xb�jN�T���-�#@,�en�(9��$�\�M�F������?��5���q�+ă���z�I��9
���]C3�x�A}:�3�!N" �*�i�,��<a�p����GDL��q��ÖFd`�����|8,�
`:������E�1|X-��Ø���í�E���-��$E�l�s�j��%�];�"���/׎�(���D����'�%�מ��P�Ղ�~��﹦1#ӝ�JWn�{Eɩ�
/`��h^�X,��v����=gT/n%vjB�j��q����kO��/�ע�D�����]���"%��x��.Fw�$��p��QA$�8l���V�8k���E�,�b��qP�����E��K���T�l��̏�?�=���Dz���E�tV��9�X\�!����o���Hr�*%	`\�/ss��K�҉�G)�^��Iltl}q����ۥ2�> ����� P�]C�s��3�ތ�A��k���y�|F��|�ѧ� K�@��E���}��s��Nd$#����I�*�ԛ�x�޸c��wJNf��
E1��%�l����SE�ǆ�C|rEu���I���yA-Ē���� &�1��YZ��,2��/&��٦?QS._G�5&��K�����
f����kE��0~��8�^B�)>zS�`X��1niӦ��c�$w�̎5y�@��A��g��z�y�G��;��7�9���]�'��󢴮Ȟ��w�di{�P�b9��r�v�Y| ���ʘE%��i5q�o���C<���ν��b�i���W(��JWV,i���ׅ7fI�ŕ�6�ZPb��0X�Ռ�u<v�-�7aX-�GE��I�b�ȋY��oͻ�g�+\�:__�R�ͽ�#;��O� %���1d���3y�)��N�~;
tx�iFgO�_����b���E)��!�4w��
/d㝍<)*=%����쬍�6��~��G�6���i�\�ӡk2�dp�j�X�M��K��\��h�i��d���ˤm�J�6����=��IR��A�T0jL�]wWW�0���'i+1wnU���%.��݃E)ǽ6�!G��uR2���j�2�w:����(�u)>�uC��<�jB8P^Oe����m��Hr�v~�[�O�_�2�ũ�,Y{����z�ҋ�>x���H�jg,�G����M�S4�f�ㄉG��)�*���Zʂ�,zϼ�oZ�EP5eN$<�{�4ی��&E�mm�7��+�7������@��ģ�)v�$�2��?�u;�Dj(S:%��2�Wl-�p[)m]g��U��w�Q&�G�#W�)�d {�}s2���'�µ4_���i��k4C����lc��ix�Y�G�"�h"/BuK��(Y�,�㑀c,,^X�f�-ܡ�66K�+�/���S R�yk!�ygm�\���yak� k\2)"��MV���x��������k��=Zp�>e#�]F/������9���/�K�ۙ��@���.j�%;�&FI�3�\��Zn����ϰ��wi���&dK.���׸B�h
��m�|y(�Y���+���ԑrU��qS��8�����y����ű��Ѝ]�ȇ1c�<���3�������ꂽ����{�17���/K����e-_�e���9�<8�)my��%v����/~�����g�)d��b[�����z�;PZ��-�G?��4����b��! z}�ײՆ�i=��`����3Q<�PTa��`һ��I���:ΰ �WS��Z?��>��/�e�NWis[��M�OP��Ӌ�I�݂0�5/�0��|n�[�����Y>�?�r�8Y�[w⯛��DU�&�e�A@��w,�paM�P!M�c��D�B�t�H)w�GةT�zZ��^1\-ǖ���^e�C�%8�9�u|����^ŪV]j�1y5�>�22�m+H�SW0Į�0���j�+(~���{�uBB6���K��g=��	��st��%=�w2 �.��d�E��>�%�c�@a�e�Z��5�"w�R��ruәǀx��O:�'?�V��P{64Y<��3D�#�^�	;kP���h��x~�B}���f7��,�ڴ�*.r�ҋ�.��G6o��x���d6zN����n��ٕ���C,4�[x"���ᲁtYD8xtk��v�B���~�~�s���>�|�$��N�c���,a���"ʊ�xD�����)oa�U�Ʊ��򍟖N�mz�ʤ�W���0�W��j�↴�\ư��|,Gʀ�D�l/y��#;����3��ON��%��%��^3jR)�)�L�������zZY._83���I�%@qd������'m�����	Qq�����oH��7o�i�mFǄ����v��	Fj�[�8$�X�}DNR�7��5Ӧ)����2�א{d1�#|Gι��I8P�U?g	g3;�U���#Vw�D�ҾѮ�����X=ff�v��?:�BW}Ij���MG���/���D,x�{b�&ӥ�h�<}�~t�a< �#G3^����s!��U���/�'��k%V���N���5��:�]u�� �")̈6!&��o�G�E��	����}Zp�h��erӀ,����.�����]R'�Hll�o+����<$ �ѹp��3�
EMY�%�OГ�	��R}77��x	�n_Mr�%�ƹ�<mcS�(��O�6NW,�^����v�0���c)K��p���Y3Z�e��d��s�}�QT<~\�]r4���|�hs6ɾe�����-� KJ��"lޚ��6B-L#�Yl�����ߥWY	J�R
Yc�v���f��[�	���O�O��8}�/޵A �,�Jc��|1��% e�U��o����2�A��j���$Е{��!�#"��C#�}>
	\C�P3y=�2�m��*�ܐ�����Z�_�g�T%WTo�~B��A�u_�/\�(�
dcP�a��ǼTV����\u�;��C�F3���|��ʡ잋�	��8 cS�%H�F2�R����X��Kj���fv��4oT�g�,'�>�u��!شtFV���������\�XZG���c�HI"���$]��DިΗ�	������^��&��OX]y�ꮳ�y�����]�����{i6���� b�K팽�if����޴�}�wS��t��!��1�	a".堀*�G�A�
|������J��"n�7�9���Y��|g|� �$����(|נ��x��9p��P�����z��]��R1e)����pY����5<zd��?�l��f+=�y3�kJs	H�{��:�{�7�����&��7�H~�V�CԲF�u������U���X6m�m���,�2LǮ@�ڽ$Q��59�Je���ޝ ���4�3n��_\��[�.�;I��Č��*Z8�*����"�R*O�RP���
�= ��`��4���U!Cb���T0��2n�p+���2O�dɕH *�v�O���$J������2�۟��b��_�����0tr
��ި֭C�{����$aO�f�`��ż��I��k���65Q����thD呟�h����x���4S�,O��[���\�̆�;�/��M
3�06@�섌�Ыfy(�����P'�Vuɀ��H@S�gdNDY�z�lS���.�b R�Y>60.U1`{��9��7&�2?M�0��S�.V�O(��)�T��{(��G����w�PX]'��^�Nf[���zUmf=�	.�cu)������fek\ �+1�$�L"i�%Z�U7"��i9b%��I��������jَ�֔6���"�ל��3_sto��zLO�֘�]z~&����?o�q��V�h�TgRI;�ק���x��kxI14k�,���Z��ġ��1�j������s��q(������{���� 2"�\bP�`�K�rh���\�u�c�M�P�-����E��|¤�W;Qr�@�X_��_����B`���H���h��NV��i��%�G>|�z/�5Y��� f`/֡��6�����٦���~�w5��K�G�IO�۪��ɝZ���+YF7�,%>K���"�b���]��-"�W]�:u��ex��8�
���C�s��T�qQ��j1��g�%Э̦�m3��=ȡ����@�ͯ|uO�"1�1s|�����'���50˞x<�<��I|qD\,f�M�7�>@�(�Es�:�.$�����5��,T��)�y���v�E�:O�o�R�_��1���3#�<"1F���_��e�?B�RS��܎0��^��U�U˵a���k�a��F@����~�� l=����eR|�����2^t���ɟ�HQOպ�K��XV������0����c��{	Q���Ϣ�lvnv �eE�V���ű^��4'�̌��u�2�$��{���w��/�ܣ���p������{Z�KbWz��Pi0:l�1ru":Ux��W+��K*I��\�C�S�KP[��79'��ZJ��kws'vo�	����JP��ǻJT�JP�������c�	ڂ��KI��g3BB���g�0�d��wУ�Nǌdg�St�˞���Z���p�J��xw���(�9�W2��l}%R:��-f`�ʘ)�J�,E7ή��h��>�Nb��G��N:C΁/*�7~(��}�~��3e>A�b��R�9l�����X�5��D<^��h���PG"-(О��W�	��:���_�S�^k�g�Ť1XV%}%r������5A��4eLM�kb��-1��j`ӳ/�Q?�ΐ:;6�Vd ���u�`ʫ�3�4��>B��Y����^i�%����(��T�++�؎�!�٬Q�7`yH~>W��=�"�FqO��Q�}H��.�D�l��.f���Ƀ��ba��-m�w���r_Ϳ��sTط ZN��p �f9N"��K}���G����Lek���Ȓ�T������{�jDA�+L��z�����bE�;U0��1X0U?��;W'��d(����h�M�k���%;9�q�jI�2�����r��RCR�F�V�k�)�<t�K��m�P�T����
����������k#�NHb]�^o�0N\`��A�k'��o���V��	�OX���rk!�]L^Iٌ�o^����-*�M�4�d��A*���4�om
��I�m�;�Z�A���c�r��V�;��L2�����:TA��3�Y�=T�az���v ,M-6���%�!����I� �jN���1��Qt2�]�ۺ'�k�����x{�W�Em�&��Jg�I}f��8���j�ճ�pt�!��BN���Kjh(���7��U�g�N=�g��v��2p�lz��ނ9�=��^���N��{zFo��b�y{���^�[*�%���+ԋkYڭ?�^BZ7r��$� �m�c��t����M�|��c,�B��}�/��n����vR��;Z<��n��I �F�,�;ٖ2u}�"���Tf��H|v�%�?��@�֞� v���i� ���z\�O|ǜ/Q����V�ER�p�L���m���,��k���� sf�e/x�`;�{<��\J����¹ѐ�*����{S��ƒ���s�	2K�����rQ���02�@r�E�f�.�洵�N�b��}LE���}h���m�`���\r)��S$��!Z؊����`����n�/�ǲ>fG��:��̓lc|�i ��ie�ڌy�@l��-��}��\���<800dŜ;�	Psp��:�8w[�Vv[w{�ޚ�է�`}��L��.��i;�1-����lC�B����G�:Ϯ�9��eD������&&�߾������|F%�]�Q�� �Œ��x�<3��C���Ƿ�P��b�5��f�%�Iy(�G��Ʉ�Nn�ɢݬvA֮g~	t�Q��_�a:�@)ȐsiT�@e�[0�˿�֔���Ѫ\�N�ʈ�-�)�g�&��#����z��89d�=J;/H�b�lk8�ۃM�?���$�ʧ�F�^[E�g�f'��t\W1P?�כL.�M��]-������J��4:�ET��^�^��-2l�;z��t���C�mj�8w-0�����A#R�_	��I��E�9�9�:'\������n�=��2j_gY!�ю��7_��I1�;��k���Δ�$�3�?eV��4�ʭ��2��X_��J�$-e��6=�ɻ�b$!��Fy�1����R����	ֺN���b1Ͷ�?w���+cb�jn�t4�`Nl�tJ%�hOJH�*�������2���8o�M��}�Y(�׷XTf�apA&8:��]#O2AYG_sW���q�/l�:P�`�������,���k���
�.a�Gn̶[E[���QHv.��i��P0���B�N������@�*{�0ҬxkuL~�SϽ{%�?���C�p`,����[�qi��}|ȜEA�
Uj���m�cR�R�{8�d�%G�<�.Q�v�iDڽ���:���](7�F|ߴ��C��e�R�B\)�oS�� �<�]��N�hZ�3+g��y7�
�u�y�/��M�`"G�Vf�U^s��N�Y�l>#�C���^q=� �D�W��8�O��O�b��' �μ���~���
ӟ�ں��FV%�Q /�&Z��x�;�G�AW52��[�*�at�C�ld��_�rd�-��o$�̏w{�0{�Lc'��Ĩ0�T������_��4��=�H��;��3�/�=v9B���c��$�~��y��� �R�[5v�w������k��k�4a^_��NS �fo�T3>�ؑ�30�[�^'����u����|��˻�Q�*�j[��G$�={O�\e9NCI1��L&���L<s�	�>�i���Y�y�����^���qO�<?�㊽Ј���Z�K�<�L���4��i��ct��ˈ^b��즨[�
������?�X��(���8)TH��*9'����*�R_�hTN\�'c�綟�g��+H�(�jQ2G����rT
��/��E%�u�h���'��]�`�!<�����.�Y5�R>���?�ݵpQ�;��}Yc��c�%��s���O(^�M��`�c&I
�'��F�p�s�u�y.mn���sZy�) &�r�ذn<���7@�9 �Q$݁/�Z)㾠������+�>�-�2�c^�!��b�����oEK�
�~+�zmUOeQ�Z�%{ l�t���������P5�ٳ���^�a�:k��y>J�h�):����7N�PX��]�v'?_�<.�!���ɚ������0ᣮ�c�H!j���X���W�����HR���_�~B{��%�>��Q�K��@Z���K|�Oe��V���r����~g�=��ˌgi%6i�G�L{��k�?�2�!��齩��
lT^�_���XSJ��s�R�Q�Gb�s��N�U���J88�=CD?'�2~�-�}���aA$�9Ž
/!���M�X��Ѱ�~HP�7��d�n�t�_�����-n�!�����ڲ���Z�AzY�jEl�p�3�&��2\��7�C�W艐��p�
� ��V���%�B�0�[�����<+'��-��4��<�O)
b�K%:����]E�ω�����~Fx6^Ҝ2��R�Ϝ���8�QŜ9a|I�}�wE�u:�N;0���Aa�$T��t'�q�^cC ��K'���L�����Q�")��R%`����[��m�ce�1��6����z�)�R�u-V�Ɨ��p,H�TʘuA�gK\����!P�y��6�\��1�|�l��i�أdz1v��� �Zun��ߩ��^���tݦ��S���:#��C)�k^�1�鲢�R$��.���
����s�FĀ]귡_��f3��_��m	��^(?��$�>����q%�K����fPU⮭�5�\Y®�cN������Y��`�y�\�C3��@w:�*dx�@��W̧Ovq��S�2��@�tQ*����<�����rE8��9[R�ٖ�L`�p���}F��+���Zޠ�.��Y�w9����F-NE����Ζ��0�|�`�r�/��͵ԕ��	(W��6;����e���a���~7r�X�z.���g睺tS\��� Ů���SpL���i���܆���g8ep4' lE{�:�������K3p_jn=u	k�v����̶�`~�n��I�d���g/m1���Gbΰ��\?_��V���ŵ�(l�X�0�ꎍ����v�{�Vz�v�B��	����b G���)/p|��M�H��"?�C|���퓧�g���V�p����B��:qA��@Rx��=⌶�r�~��	���7���}��~����`�PV}��$0#A����\ ��bB�H��{u�B��Ac4�>����
k����Ϙ�����r,\�o��"X�_]�Lϒo\aZ�6�����:���SX��Rزˈ���MD|����: �=UΜ:%�Og?��U<Ίo�T���Ж��X1�P�o����0`�l-��N��?[��:,Q��qQ=�OO�y���$�焝��Hѭyq��VЅ���]��<f+o#�1 �w�~��\澻�N�-"����>��)dWga5���]v����u���u�&���dM��E1���F��>��/Ќ-x�����]�H����K)�+ʐ��(��6�̞F)�u^��,�Ankxg�h�Av��Rb�j������B�>V�j��d.F�Z2w���'�ڊ���,���QS�8����AΡ}˞.
3�%	�^��y-P�~`'��n/�X����6�C�q����k��㳒�Y)���C��P���9D�
��� ��j�T�90^��'IaY�i�b�!�e[:�n�e�+U��>$o���؆6$�g��J��{DFL;���/��r@XUx�eq���O:
�����-�§�`�\Y��)ץ�*����@u���h��J��x�E�Vj��=E�^�;����wf�B¶�>�����/�F���A2,����b�_]����i��$_5Kx�#�p�q���a$io����I�A5=D:���to��u�%*a��\H)�o�C�4�����7`�H��R�陑�'xmZv�I�q��W��@���n��H�{�&�"��/�z��ɢ
#t���id9��#V��F;�ɇ7$�eu3� f�J�!�L
�u����{���S}�F��ks)Mb6�2��0K�H�}_*��a�C�'���ɒ<JA\ac� ����N�\I�`�t#x�Z��Q���4#�z(�b�V���^���3hT�Ho���^3��9������7�+fO�s�2;�_�{��A`����i�Y��U��$���4WJ��!��85��N7=)V=.T�r�n�x�(i���U|��Q��ԭ��ф�W��%/�w�9��z���97��	'�ΜtRԋWA�����q<XJC�[��4f�\��,���S����W 72S�B�	�&C��@�C]�X��Y�e!���h^2n�+i.0�}�" ����r' �m_D��h�(r��	$_0�����k0?�*�ї�Ve31f���*هQ�ȀmY��՝�=���a@�ƚ��1�	�dM���%�����R݂�\.�wNɃ��Zҿ$�]����fV���`�M `�����tνUW�]����x	}4*U~�>�E�j��Į��{dB��#����qҢ����<2�>��%���j�*�$�� 9��'�6y`7����	M������a���W=l%/�a>Vk 	�W��/Yk���"��J�9�\�<�3�=��W��$�!`+E=�OII^h���%+�����n,>~1�|�&�
�����T!��Ѹ�{��qb�f�m3������إ��,�z&�f�M�0h���W���VX|k�T;���nYUP!��B��C��
ޮ;�����$���X�w���ݢs�9v�4rmz���O�ؖn���7�!9	oԮ��Ɨ�$�(�X܌�U8�)M#��z�K�^������i���gCd CO_׶���ߦ�����hk���:�\==���׆&G��	x�p��2�u-}P�u�����]W�w���M�k�܇��lbY$�>9��8�=�_$�N��-K=��mXk�wl3%&����C�F�a� s�p�+���7�)�ɛ��n�eD����]Un5&w�w��i�E'i���[e`�ݾ<�u�H�O�ev@�O�����H�S��=7�lӐD�&�́�h2r����%I�����(0H�~:�WA�n�n֢'
A\���DZ�1���Lz��w��]�{�:]	N|��ӎ����
`��,5�R��A0Rc��.�O�b�{B��́�G�A��2N9!��QO���2�����T��>@���W�Q�c���T�1p�z��>C��y	�t��0}3z��;��l�x78�u��!�Z�Wi����P"�j�ن���Ȥ��\���� z%�B7�T{ޒ����o��'���(<?	.���8��O(s7W!Vَ�̌/v$��[��f�~�{��'�7y#%�e�\1���:��B�Ģi����(v��6��QzcE��pj�������MCR4�y�,���A%�&}5;����5 s=�&���-(�G������#ס8��U�l��b���ժ~B#z��T�w󌞛��G��#b,�Ă^h�ﲱ��(|��7��9t��Tl��"]O�����~��?�����.\?\����<�a&��A%2��Dh�X�p";�|��{LUolp��y�n�)Єo��f�A=�脄ڴ��2��<�M�QS$�e���U���Y�S���v pBdM�{���uW��?�:���Q��&���u�m��.�;Ȱe�*�3��F�_��������@� ��L5Z�����U���]sg1 �^m%6:n3��u���n 9B|+��������p��(���i1�W:OiǦ�������v"n]]>b��/���k�L����8�p�^�����m�EE\-_��Jr�_�B��WO��t���ɰ�����=V�8�:d�� e���6J9ʱ��b?):�G����ˡ( �8�>X^N��階�O�@D՞r�Sp���Uw����w��ӻ�����gr@n��B�̩�aދڮ(i}��!WÍZ�4$O�m��#%���@�/[+&%=o�	[�@<��(
J  �Nw�?\��-�����=(j�߶��x|[��@�K�Jo�l�
d~O���M�4�l�\mx��H��*ŹZ�-M���k�3RW�G�2�ַH�Ww��T�xu�Ğ8<�R��_j��ٸ�W�6�a�Q�E�a������wm��3R�dD+�*�QM�l���2�0/��6H���rǧ&r�J-8�p� ��b��F��]s��m�#��/�@B�y��b��&>��l�M��k�c�r?���|8�l�K@��s�]t���ڟ]
q5>��=I+�f".��)����*
���3�����V������{�K�@혥I�Jb�����&���d^K��to�� q9bWF֤��#B�r�O��j��!��Zb���V����0(�Sӡ&|V�b]%	9R�y���6��𣑎�c���*�rO���N���}��㉯�BQ��͔�]Es#C0*8�b��������Ruo��dgaU�TE�_d�қ#�g�\<>���&x�\���U���ɗN��������=��ڍ��I"޸�y�|,b�9�rb�b����A��.~5���E�FV�v�-�S&5��5ĺ���n�ڙ,{	��-t�I<ێ��zu��y�Ґ�@Mc�A�x=2����q��a�'y��	�������		��� E$�=
��w��Nk�|U�MV.�E>�R����K�ޮZv$&�S���ߘf��'wT@��?�B�gNi K���[i)��O=�ʥ���爥�ވf4�x�n͸=L�FK�'�WM9���k{?��0���j����G��@D�KU�j 3o3��I"d�F}	�V~η�ц�i�_�ΟUw	PJ94�It�4���l�����q��O̵Y�u�?'���&JƧ�{��C�2bޚ��J |BIרrO)���S<��J�4Xa+x7h�7������1���G����	MxGSԲ��l.f���RcO��wjɸ��}!"%��&0h'���{*��҆ �����>R��ɽ�ş�/ 9�*����Ln��jU�;��^׬Y��+��N	�CxO �8����)0>���y�L�l4B@b9i�� ך���"�w�^�'���_���3�l���_�W�)2H�^XVm����k��)U5�k/�f]�rCa���gה�9��!�Ko�tV��7*WfY����g�6�Mҗu�	�]V�����GF]ɻ	*���˽�U��=�]�	/A�<$8��z�ߟQ���)#A������4�Ea'UK��B0��V���ގFR�0��C��/ v��{kn��K]�Y˚�5���lD͛�Tb��>��ބ��U v^K������x9V���Uo=�3 6����6Al���w�|�u^b��L-���~��5�w�K�"p����۷YZ��b�����1�>���z�Jl�����ja�%�J�9�V���j��&==D<�>�;��NF��<�8(H���'��s�It���'F�qD+�Dj���\�y{Gf���Nm
f�ָ�y^�b��[���f��3��e����-�w ���1�z����빍y�I��mr�~/\�Ho{�kM����ƍ���X�5������X��"ѡ��U�}cg�,��~KY�:���sV��5����R	l���$�r���8"��`s�~o�N��\;T҆��O/2�~S�&�Ŕ9e��T�~�%z���(�.IU+�;��o��,��0X�ޮ)G�Aݸ���e��Z�`�����=�;�ڳH;n��O7�j���*�>J/u����$|��`oQKU5�p��4"�/�\g|��r=�vo��߈���UL�1Q����6)��é6"	8)�	%�=r-����G�+�ǃaY�HI*�?mV3៫C��4o�-J���Hg��)Nk0�����v">�"��Tv9 �U�R�n�r�ۧ�����f�h#�I'E����-�8K�^���s^w�)���xP�/-Nڋ���{�BD��r��g��7���Y��K4� %\�����֦R������zt�Bg���)cS~U�+]�.|$��O�	�N�`Rf~�w�bW��v�
Gg���X9�!nN%!�~�t�qp"�Q�`��f�H���:Ɍ>��+m�6f\�8���Ѧ�����A�� �zn D�����$&{%�`ꨏ���2�2�U�ȷN|fKX$W�k�"F㸹j?�l�����gUy^���D��ӻ����Y8֫�(��7�O���[ؿ\�/%Q���Q؀�A��p�o�,��<�~kb3����O���a��ܔ��C#�(�4�YTv���Y�
UiAڬ�B�a�n�o�A�tl����ر�4�|I$��b�����G��D��sjK5h)�b��w�43�3��#��2����ED�Z�XT�P\�R�I�>7l9��ަ�Ǚ�����/Z �vK��Ա��M�>ğY�2>����'@zw�tO�i��+"��ݽ�,Ċ5�īJ����Ѧ�rf+�ʟy����(n̇����-���U	�'cL�
��E��.�-J�t�i���Z�����{�g�p���S?uOI����=ِ�\��� ; >�Nv����&�5SC�� �� ��l��l����nD[E'���wj<q�C�JA��l�'���ē���x��6Q`�O(�y����r\�r,��	�>^�1
�G4͂J۞YtRn��
MV�[�+����Qr7�����v���H��J��4�C�>z�@v�\֩�a�q@�1ci�Ǩ1��Ӣg���WcS�d����!���;#0�1�C���{����o�θ��'���B;b�|fN^�->f��_�Gۑ ��i��0�
2Jћ�
�� �E�X�\����X(
ˠ�a�s�D��ĢӒ��E�G��$j�����mBֿ�آoaJ�y��մm��>f�����5�}��d�ĉ[���{)ܞ�*�8M�z��B�+����i�tɛ��_�\Q�'|��LWw<;���d&�gn"����j\A��+ ΀�T��,�_�w9u=Aca��!E��+n3�1�s�E���x'�n��W8 "��2#?�咞����81.�$¼i�/EN&]�p��������!�Z��H�=�fG�!�ן��������L��Rrlu��s`hp�E��h7뭬��͊��жKƺK�[�sʛ�ʇ�d��~9�������:��̼���	K��� �[=�ے�a�G���۶�����YQ���A��=��M݈
W��5���UJZ�j�D�`>�x9�JU1�ɵ�nȤp��P���0������S�����H�ן	�sgq���/��=HA��:$�#+/UrŜN�]��=��[�R�h���{��
�f�Z��t�?�ҽ�53-��z�ȩ&�KM��(�K����A�	p3�	f�v\wGy(}���+��?^с��l��p�o6�op1H{n��M���Xp9�ɟI�ܙ�Ί8�o#x� �z:\g�x�g�,�cό���%�i�.��� mE&Jv�쀯��у�5�����1���z)�Ƒ�6/�O�����ߒ@��cF'�/�I������:%d��6aauJ�Hi3�V���1�����fE��~���b��=O�~����v����z�n�!�б'������Q{��cu�<�\�u��e�|��n��T�B�z슛k:�A�^��2�S7�Z�J���S�իB�|Ξ�����6Z�2/�b���^ُ�f�?<!
��L��3���j�Ct�Hׇ��5�1�e`�a>!��xm��H�&0 c0�K.�GC��7�Z�G�D�`y9D�XE��A0�� ������%Ѡ�l��S��錗�z�<wqӯ?�8���2��f�_o)ʷ ,�b>{�$T划ۀ7T4��)j��B�59�.�>\�TW ���!ɷ�������.KZ	�uo��-0@��mLzy�Af����N;B�<����	��nP���S����b�b�[�n���/�Q�"v�5���`	�H_����u�Rt`n.|�v��i��x\��vDT��R���m�ۏ���������ɹ�^��	��*���M�T3�􏍸PF��A���B4,���tZ5X��?zn9$X&�u��W膞e�Vɂ#�C�Y3�3M���$�J�$l���۫.��>AӞ�P[�bC�ߨ&=i��ZHF����qh����^�^�%Ÿ��"���E�|�~8oѹո�������Ce����|�9�v���%�(%|wv����Q�m��î�Q�O�@-4Xj��k��
�a�X3�c��G�*ü��d�о0���J�6*�aw���7c�k0s�mWUw4�1ӱz5�i!��N����}�ތ���Yԥ$ɾ	S��2a1��*#��J���|��T�є%�B)gU$#[�F��z�: b���W��p6o�Z�=ġ���m�