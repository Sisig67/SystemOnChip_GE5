��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%����!�rr/I���b2}���Vpiv�o ��g��(qα-X��$�qڂ�]Ub��?෬�H����|�t�Vo��<�X��{�NookK"4v�
}B�ݮ*ԯ����o�"꡼����Q�_"̲�`Ѕ�-R��}��v��������� ��Nah
�=Ѝ��oz���^������I�&�Q׷���>��W�@��H��b�:�R�CK���;cOU�M���6�cu�W���hO�{}N�E��?��P�'�_�C�XO2��(��1?Ï��`./�({�mP�(<�����4Y2�����ܖK`�gnb(
�G<��HP��޴�PL!r����]���o�L�vDt)�gK������mp���Ami���!����@Bs �0k���`�|��q�iv�v� �l�Z1#�;bG�ȋ��w<���Zg�9�x�Fh�uP|�sGF���j�wM.]��e۪>J���v5i�b0��P*=>��y��vL|?!��h5iW��l��ʮ��#���!����rS�^��.*b-�����^2xݙ=�	Y�8�B�>�~9s���{hɾ��h����K Iݳsmx �΅f��`kz�����p�ٹ�B�Fó��&>�
,,��n%�gCΜ	��x!��r�6m��=�UD8q<����t���#�#�Ln������h��9k'�L(������4�Oz�LSwLͦ� �3р�n�wd�[aMǃ��jW��,���F]V��H����!--B�2��(<�ނF�[ny<B��$T.C��Ɔ˸��[;���EP�Q��2�}��;��1&\�[:KO�e�Xt���!!�6�D��/��F�X�Px3�m�v�!�o9.$Z(�D� �F����"���.��{����X���G?-�{���^3'�&����_�==�3��C��Yu���D��:g���U�q�9ߡf/v�@�HGCej����vN=�Y���O��̓�y�s],���K��=C� !Q Ld�+ɇ"��Ż���b�@���vl���-WQ��:z���a�[ID����dL��.ԍ��FB�dZi�0s�X�E���	
���� ��L�~�/Z?��I���{"�h�L������=V[;U�|������]���'�+�vL�/�9G���)�4�BJ���Q'J�SP��}К��'R6�F�����6B�r2~6���?P�P!u}z=� t������^,�@��2�u$ى	���wzG2�^�ĺ��ن����æ�1�!� �,�Tld�Gw��p7"��]�h�G��0��`
��d�.Rm�icӺ���(NW5�����I)g4�>�
����Jˮ\�*{�jQ����d�y�`�9]1���T2Q���H�+[��LL�O�-.���8O���q�e*<,���Hj�c����rc���;��;��
���ۿ��`ِ�S�"�ѽ��A�!1������;m�[ɽco���J�a����se���wܛ�����cD�G�����'�����g�!�d5.nu�xG��bK�4ǻ�J�'�A�:�3�[��
�8���4&��r�ҖB���5�|������Jg*��1�I�m&D��J�wDen��_�x���v���D���kn��󱺺�=Iƒ%5W?$yBw)h�"��3ZL|#𫑣����F��]�US�h+�1�&֐lk��UW�B���,@��/8���ۙ{�����>ރ<��q�Nѐ�?���Ao���+6��T]Pj�et-��B�Q2�vQ���W�j�L�G������EDn���[H���G��T�5������� ���b'ۦ`�R5ZĨ�,�3[;��֠��Z�����dQVܙ��P]��9�Q	����PZ[#Q@��Z`�N^�d��VM
��w.h��6�l�(�6��ĥ2����z'��c����ٿ_~������E�b�9�k��t?T����J�\k}�����^��s"7y�l���ΤV?�����)��z�c"�g����.^U�T��gy
L�Δ��4��-�-��G�'S��yV�^�\HkQ
�M����=Ƽ��G3(�y"z%���~P���zo�=ѭ��@5�q�1��� ���L�e��-h������צ�]4*����1��bsi}r���d�v�m��ؙ��a>�R��?�6�L����¼^�aT#�3����9�N� {�'���t��f�r�L��J:~G8�k	���:����2=�i�Oo��Af��\����k�n�V� T��	0`��Ǯ%V�n-���[�\����J����
�2|��������HA&�<�v�0��º�a"�V�Y!�Z��L��r��Yw\S~���<+�h���m�o�2�֨ۦ�,)�z�/Z��� �K;��p�a}�0�u9lU��VU1�m�u����e,��[Q=\S9R������e&`k�N!Fg�)����R=[Jx7��ж�a^ypy��3q��"F'2V�_[���_#��>�O������).@g"+|��V��bN~������@U��`���.b$�E��4�g��%%��YH�*�n�����^�.���M����� "�(@1���3D���i|����#��g�45z&x�pF�b'�`��@#�U෵�jG�Y6��,J�5���gyaT\��#h�ت�f���ﻔ_>��p��s12؛zUTBE��S�s�O��S�m�C�zl�ۃ`�A�.9�K���}�i��+cA�)fdec�Ͷ�+�i���z�o�vʪ�u+��9d1�Ҟ�@O��ֶZ�����<.�!����w>�Ȳ��̿*	��9EI�=U9�݀D���R0"��z�=b�,(��B�C']�+
'٦,��x�䌁<�;@pl��"���g/ZT�!	O�,��Yt�4�zM�������<O��1�?Zz��ff-h(�G�.�ڵ�vO�Lʕ	����0g�G�V"[�̋���B��{�]Fc�|�^�6!7�8�rq�c���#�eB�i�|�<��w���3@�u��gM��Z�=�3I~��DB��`�r��2*7;�+@p��-Y�my�f����)@�`�Jj8����4��SwG^�vX8տr�6�#��c�Ʊ��G��t,&��]P����Y�|��'|+R�2�yw�	� ���d���n|zpd+K�I�8x�HQ����5��ZȳJ��� `�!�u8��3���A����C; �ծ��	W�#�]��*�`��H���{��`Y�u����	��֋FUBV�+ܙV�M��wC�d@�/����09d��������˴�C'���Әy�3{?9}�_ސ[��,A���:�,'�4j��{�
|��	��N�L�JP��X�����Jg�C�o����I���]Q��
ةz������4
���`%�Hղޙ�]j5�H��qվ��%ƢB��Q����ǿ���;�=�����-=��5�_u�+@�ӫȐ�R����Y�)9O�(��Hʡ+�
R�&bw�����c;>u��wz�hK �Y��J��������u��GdQtn�)mVc
іh۱����L����_U����/3��
����&)ъ�IF��C�ؚ�=�&:=qf3�s4�����R�'F����;����i2�!&��O\�mq>�6�V�͐u�ja�E8�X�D���\�<��y&�*
�2)o�o�W}Q����2a��f�*�
��E���Z�����)�$"L���2 6�P��#��g�}�%�;��rv��%P��>��Ax.�O��<WR�iz��l���T<OnY���W"NxbM9(��XYX���U�b�Ś���53�W孓(<�W밞NF���*��p@uj��E]. fw�J	9l�8�^	D�
!8~���7��C��M.a�'xhp[� � v=���|s�>x�����<��l�J�;2MX>�de��PY p��o��˳��A�W�#��I�(��"�4,��<��H�"��S{�7��1'C#��T'�Ǧ�s�g�I��\ Qr�u�Sķ�	�me�<6i�]Ī�^���ϖ��g�cr��όO二K����cZݖ�[�5�V5��5���4ф"x�sL��o������xT��DrWC؂Z��������+�܁@iZ�!����5G#?:ub)8�X��CVg�:����mо2.�/����ж\����D�D Ml���7���!����Z�N����ךMj]3�:?Ҧ�Ij��ؖ�YoX��L_}����("/��Լ!PD�~I�+n�N-v��]���ׇ}��K��;3Wۈ�� WX���B�J����.6W	P��/_�bd���O�t����A��]=U}���$�e��3~�=�=�,1��n�zPn1�Q>ő�m�A r�솙N?�o��2�QIA+^���:\��9+�a)qE��'$8=�� ��G�Fw݆�8��-[�wq�%�1>4��!���<P9iI#3�#��S��ʥ�����g���|����淏�zEm& O�Dp)!B�w��� ���#98��oA�-�����Ά��Ry��P��8_��#�=ݕ�3�V�)0�|�������o:̋�!���,�P�M���؜e}W�~�N�9X�s���V�j��	�:,m��\�!�:Z�JB�r+l�N�QP�@£��8]��G[Lp���r�����/9�-Xf����G�9��h�X�l�B´:��D�žt�y��Xђ��_�K�߇<f�Dn*\<�	�H4l���y�"/��g��.5&$�� =.`-�7��i�S�B��y�1���*O��x_Q�\ 1������j؉d0�7�ŗ{"w�e+W{��$��t��.�x�����{o	٨|@I-�~٤'�_q��Pz�(��_5RX`q������7⫬��b���K�;��*�hJGr�����5���U�gne+"��/���Qq�0��i���Ú�YQ���q����=��s�<J>��5q��ze3���&&N`��K
X�j��ԓ\K	��[�}�u�~_Q%�5����O������� t�0�z�픒��o
"�h���q��X���[�������}Ӱ�߸�RA=�b�2����ރ��s�X���Twg�:�sS����U���ٱl���-�;K_�zݓ�7:{��݆��9}����j|�0�&|Z�zȁ�u9$���訯#Oh�l����C� ��x1:jUZ��S�KC����)��G��H���X���s�7F/���Txa3����C��Ds�p��+
_T�Β�E$"�S��,hb��\I�TlUz��@��������`Q"ȇ�2��}�x��o���q��d͢�~_;�%�ۘ�Έ�_���lO��X
��9�M	���<X��-{�'E�)�v���h-�(hjt��ѱ6�/K���ͦ�d؍U��N���k���c�j�⡱\�Ω9C���i�;�t�ў=X���kι (�~�~��=I4�����7`pJ6����5�Z��;(y>&�&�:p˩J��3Dފ��r�򓪀����V�;�SAcd�r�u��km�a6��kն<y���Ý�G�j�W5zBQ�Ho2:O�Y�4�j���)�y
�;[�Tk�ȿ���ޱ�jӢ"���0)�`7��WLz�� �<�L{�v3/FI1�)�2�}��8rOZ㌏�f�W9=�Pg)���?$��9H�J�]\9o�n���_,�$;��\�K3j#B˄4" �Y��P�G���&���b]�1�+z����'��~������;Ɂk� bM�A������k�E�����FH*hE�=Tl��R���2���3xX@qvî�?�m��8N~oB����w��N�K�����l�ɽW��S�H9���;ޙ��yl^�JU����OH_)�g$��ۅ�MC�,9�Pw����z�q�'V���Q|t�.���5	�:���#0D�Y�B�(��%�΋�D�0f�ړ���,�'���nQ�*eh	(=�Z����N;i�C�+~�au}���YW��{ۍ 9͗/����OQ&��M� 1���oc#g��O2�F4l��F�"I]�dtIrNV�}���#`7:���CUD����P_.e�ގ=�x��?�n�`� ��L=�
m�ލrJ��f�Er�w���bk>�H����n�b̎�,�p[`���gzZ�"&��J;<e�0�轋�����XH�����P}��t��kպ��fϫi�B+�zb}$Fe��Q6�>�zfy�P����u��l�/�?�%[�F}�aG�K �yޗ��n�|�c���\g���T;���	�w���U �y����9jbۤH$k��Џ��"{a%rET�i9T�df��g]�a����z��p�͵���s'�ʽ�/v=�¦/E�zX����}����%m��$7���8�Wx�6G[L
h4�}�=�#���`�hwŝ��aԭ�>k�y
��ӻz.n��N�@�����,���'W�*�r�	��N���y 2��$2{
\U)�؉h�ҫ��|wؙ�P�**K�K�}-�$t��T�;|�m�O��M�.�00z�~��^�z�v:m͎[��?=|?s+�d���Ҋ~��Eb�[���Q�(�Ӂ�7ڏ&m/�#ߤ��k�6���!,����dC.�Yˠ�)-I�429٘
0#��a4/#��U;�ĭ��c�"B\Q�\yX�p��fXoa���@3��D�9���bB���P3Q�7�T���D���<��e���q� {�С��<��3�?K7x�
f*����}����f<�9ԤwU���	�u�7��f�,�b�������n�I��ނ�%T�0&F^9Im�P�\;�(z��Ʌ�6����ϳ(�
�M<�Qr���n���ݘѿZ*����:#S�l��-zqf*i_�*�p���
+�V\��Z����ST�W�X�
�V�;��A��%��b�����nv��%�����~)�����И;�%�����k�h"��G�,��bHβ�IB���^!��w�l+:��/�Sa66�]nl��C$�L���O���������6�RQ�Gn��7T8<){���_�*Q�4���iSH%�
_y�WtĄ䏧~�)��t��
}���u�֗0�����/�
}Fu�)�=�d|�7@[*�Љ���	����䴒*�ܼG+c�1o+J�2�ֶF�NYH8���j�ʑO\Ө�p� �}���@w��v��O:�]�u�^�n�*ώ���m`�*,����d����T $ ��kO[9��IP���8�t����b)@�M��vN^����-,�N#�10z�)v��u��ӁN�Ъ��o",%�=�)����dp���$ѧq,��l][���Ĳ{�qP���$�?���h�	�kF�Jk��	e	��т/@�.�&�Pv�*���~QI�>��������7υ�$�K�Pp�P����t���Aˠ��l {v��U@�2Q��6M	1��3�a�E����Aeʹ�e84W5_3U|��P�y�8�򀊅�*O�t����-1b��ѡs��i_lE�}�}����	|+���8k�&dE�b�i~�^]��Wx��K��u ���S�O��}_����e#�|�=$��9��@zI�O���}+��?��C�ܤ���"|�"�̉Ʊ���X��:L+����nơB�7��'8��3^��x���H�c5	[�`гγ�倭�q"g`�+p�0Zu��ta2E��3����R}k^���%��7 k��gI��)#����UmBd�E�r�c�����F��0o	�hC������`�����O)