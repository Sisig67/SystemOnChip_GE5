��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj�N���0��3�J��a
_h�\6���6��ϐ��(V.�i�f;�T����� ,$��gA��'��|3�%]h���}m8*;m����:�t�����`�i���$=$Q��K���_���п�'5i��}	�����@�d5�-x��j�Q{"����C}v���h�G����w�v ֚ۨ$	�^4��oE�����BUY$�(��˖@f���}�@웲|������Y%�n����/t��p`˕��Mny4����1�I!����?�)�XV�H�!��,g��B�3�ÕC�����K�{ZKt�4͡�J�?���2N�D4�V�<��"J�g�c,�=٫�8\������J��z�_��_�#��]���6�Z+������RJY�򡎻8G����K?0ʋ-ޔ�w�RC<j-t��/(5�%�fm�z��v��Rr��ˣ�a�t�'y���W+�pļб �w
f�4S��Ėx��kݯ�B��2�]k)���j�y��7�{�_Q�t	Z�o��@�o��!�(����&3"]{�w�2��O*d�(�����x3�K�3����S����&�cc��/߫�ud�	�	�qWkG�8WeHq��J?��wX®q����[w�S2�����H�&
$P�YG_ʅ�oK�(JI�u���ߐxA��%8�W�lV���0'��DU�%�ܝ�9@�E��U|`��{=��5�8!���Y\Ie	~!�AA��T��lx�!ftO��>�p�=�5�cw�na������g�!t%u"�n[�&�bB�Ot�tiXt(4Z��X�9�y�xGPe�^x���8�0��0��rFg�ʘ�
-��Y���Y�vWaB�Y��wYB�?�]Vf�G�V:�_�"���B%�8톮��18���[��.ڙxr��}+�J┄�7��b��uXԋl��ư-�4)�*@2��Z'=``>���ze��:��pfJ���ޜ>N�� ��9_��E���i4ߠy]/��d����zy質�7�����{�5'���>�sq��'��Jˎ�%�һ:;F�g��X�)�c�p4��agN���ӡ�F����9�.��0q���߅�
3��p�c rF��C:=���3d�!M���r��Z��Y/�nS�d��P�����)�nf���^5��Ⱄz�^K08�O��8�|���c���L�B�� p�">q�t2��2�!&�#>�`Jj���4{���_sz�1�1�Q_ړ�/�8ő�iSV%mX���"�AɁ��/�1ɚ|�c������ӿi����f�5���0 Mi#��I`�D{J���"Wr7<	��eu����`?&i��	Q�{��sCLgnՂ��}��c�1��M�N�{���`uz��.��s�98���n�<��^[#�g�'�G˓�@�*KT���A��D�m.�ͨ���/\�®��T�ؠi`�jR��	�9���m�x*�GH	�O\/�<�pv<,��>���E�,2����]�(ilF`�V�	�=b���&�� ����<�|�'HE����
	�/��e��rP���`܃ܐ}�Nܬ&�CU	��hV%���rJ�9���"ZY ���ݷ�d��WH���D+
�~NP|�̤(��V�U+YW��/��%��r/�Y����WB���o��꿴F�	s����=�-��+�T]�AZ�p3~�K)������|�ہ�
����e��8=φ�~���
x����E�$�l�P3�|4� �Ǡ�������{l�k&#Էn�4�r�_����B���b�	/ z�\ЀA��52��P,��RJ��"���SL�2h��i[���<��~g��=!��=�6w�{���$ �3�æ%Pk��vhe��E%n@s��R�] AQ���	X_�C�����x5�h6�E��Izx��!y����lE�����qi����pܧP�?ޟ���
z9�kG��g)l��KJ8���%�g��R�j"c��s(㙷'r�b����G��I�$�
G��^�b�KPh����i��2�d ��G�&���E�T�ltpc�R����:m����A�+
S\�I"����YĻJI��A3 c�@8����t������;�4OA߿����:�=p0Z٥�-@U�������k;Ǒ�>!U�%��N��]�������l>G�\X<Ո`?=����$x�̂�,UG7;)�O.Ih�B��ǋ]vł�g1�y��$ņ�P[XO�B����h)�p��ǳ�p�HF�h���Ue�s���u��k�i�lT!}�"�org�-R��?��¶NL��@|�Ɯ��T�����W-�k��iQrH\�R�;�Aț��� /, $���r�:���}¬0R=�ƴ�I�&*�ݮY�׻�<6U�Oe�\Os߻�a�.��h�4?���L-�����λ���pJkՍ�<���� �炐M@��4�-��F��>~?w¡���c?��تس��w�4�L��Q�y������,�|⪚q�8����F2zҠ6:0�����Xt$�hJR��H�e�X����C5��IY���rW֋0�s�޲؋���cTz��������}��3�Y������~˂����5|"�Q@�5�x`�ײ��W��E���f�$�r��+��H��:���B��YDW�Iɧp���@ lf4�_���R:�f6�#�J
τ��z!H�h& �Ƶ#�w �+B��&?1J�����  U�ݖ�_!m�\sV,��.g��x
:f*;���Ff��0�_,}**b�s��+�W��"3b�r1+�2K��j�oA-��/���3��9��*���3m_��4���Jbw�v*��xP�ۀ>V	'X h�Di^��Xw�8Y�8G��\z�0�	���=3Kn{I�V���dHE:
́�F��p@�/�t�/B��|=Muɪ��*��Q*!�X��UfM>H��eL�٧\O��_M��B9��XH�}�q��\��(8�ZĂj���
�i�@_v�����ٳΏ�7�]�<�r-�!X�>l�;3�H
T��Y��mk� T����:���<�ׂG��u�!��\�>'� �I���'�YI��=�-"1rd;X�p@/�0;MQş<38�)�ETnZ{�CH��Ȇ؛ы�)%�X-�\��q�4IA����&D��hd�<����yʚ ���'���%0����[�_�A\xA�_Ś��{uC]0����������R�X�F�W#�U6���{:�I�w�3z��]�Q;��������T�B�q���/��X�*�yR�-�῭��q�/���E!���ɑ~`�}V��%�ܖRp�诧�:w��9N�F���.�Pυ���`�+����+_�y����-��W��.G/�'`'K�a4IQq�OH��D}�9^A�B��`ǘ�~�4��k&�m��j����?�Z����R����Dir��<��4|bt�S�7y���\�m��̗��t��/�~�ڳ�x�5*���ɓ�c���t�8��t��oi�M�o8H�B��R�0in1u� 6�� �C�$���=C�3�����x��{@I�Û��ʯ� O�b�p������c7?.�֜`�Z�����T�0���Ğ)�T:��eC酷*vE�-��9��Ou����p/�}�f��J͑���k�Y�j@!\P!Ĥ?Xb����mԂ���*T �"�AL�-z������Ѷ�C�}��iX8����-��O#ł���L�Հ~�/�\�{�}�_�<F�}�a|�:-���	|.2�˹C���p�6���m���_&�i�h6ob �F2�]��[��+�#pmg�5�45jۜ�Q �W�>��S)�u.�P���o�@\�֏,���dZ�E8{���,˶^�a^���=�� �8(.}$_D�a���M��\j�0dOD�Tv�l������7~=G'_���s���U-�'q#�ƉZ6@
8Ŝs����|��}N�	M�Ǒ��M�F�z�ա�ԗ��%T粕�~� ��d��D��} ��|���n�*I�BQ(v�<Q�a�%��曌A�#�$HS�J�e6�C�ND'� Nq_�� Y�H�A�7ǩ���'ia�d$H��mj�"�߁��bv�O���q���-����t��ֆ�CaF�4B9	X�h�VC}���u�׹�px�����Ɇ	�<����:�L�n�/��$����ה��f�j���6eC?mh6d�)�).+&�8�G$m��;�a���{$����-u�*���F,��2�otȔK��X[��!�yf���ϧ��K9�k~-3�ȣ}ԃ$O@g]�u�zU�}�I�{�1��)5�iLo��3�T�Ł��ɲ< E��w��Lb.�"�A�{�:?�~�dG���M`K���6�\mI�=��}�V��P{��[N�^[ [/��r�z�7���4h�&��\gRZ1�FW �7 ����EŽ�&��d��~Tl0lr���[��-;�����b�E?�+&Jx<�j��s8��MGG�*F��cC�Խ���ޖ[��lr�2��d"|��+��qX������8�+� ٌ;	�5 ��W�0}*�p��#����%�ނd�qk�Uwkt�DW�.���=�B�W��>��z�na��w�Rp1<���\O0. �	���$��Q���uf���YCrJ��l.��#ݳ�|�R ���r�j���aN�t'�[��G�B;��_����<KrFx��nd��B[�s��"�d�b����7�ΰ�R�k@9�W_{���3	5T��pK]��3c��,�N�x,[�8I���$�o2b��6����p�=����ؙ�!)$Їj}�\��;k�25���+x��N�§jq�ڢ*=Z��OȈ5�o���ɿ�-_��>c�4��']E�R� yuv�fU�����45� ��{tۯ����aV��ŧ�c�<���n&"p��U�ګ_��Ч�Po��ȝ+�5�n+[�p)x�d��Z�wK��w;��q �_Sk�~(�݇灜tW���I2��9D��������rDS�)�=�D�_q�rI5����:��byZ���_���9��û��� +KC*:� [aEvm��'#N}�|rr��A� ��k����b2ָ�����L�(��XSU���_��L���C]mִ�sUU2�H��*���m���!ᗝ$fg�n$u���[�+,�����U4x:,���)�m`��B�����R\T��*�k��.�2KK���_���5
�2�4���ug��Qh�D��_<)�M��p��,�v�k�SS��ŏ�	O>#c�~'���<�z�H�c� �v��!�;���h�\e=��.��Q�=fH7u6��E��{f3���<�-�q�
]n�`4��Ga�Z�Q�M�K���_%���9�\uw.6<��o����;�M�	@z	d��p��՝������SNt\��MA���u�t�ё������_a�P��u5����n��S52K�P�uS�n�ΥǠ�#		�I��?�+�����8�oj�9�9v#����'���0�/i��V�yf� ?��f�1�:+�����]�L���J|��;�h���
�*]��O=�`A�㰍�u��:��?��lR|�u6
�5�P�jWc���/h,����I��mH r�D�7�c@���׊�{ 9�I1���ؑ6�y����9���A��ix4�(%��"*��ӱ��f������&=�����PQ�ʹ�*%�Xo\8�]tOTmaÁi1����O�{s�Ց�z�}!�O�d�������a��d^B۝+��do�1j2�hB��㴔��"��t���!��?�{O�n2�#���2�����ZC��5r���_����ÏƤ���������9�{8�"�;e�u��\��9<�z���0�O):nd�$�v�����x�ʲ�
��ih��i�N��D�� l
���̍�����?��+��WG�5�޴XO���͝��m���r�Ö��f�����"��K󺐇t����%����3��a��{�}[-�~�8��y*>�:�XĘK�R��nU���4��N���]i!aU0�łu1Z�в<����,D֔T�l㍭��q���m�-=�y�T��#nr��4�s�_�ڥzŘ*����Lk�ߩAbWX36���0�0'�ux�:�N�&��j�_��yZVu-�u����uF'��Y�������\@YP=p?���)q��D�@(�Z=E�X�J��戩HonQ���K%��dP����u�>
��se������}}Ġ��o֗�D�Mkoӑ�f-)��{�"
�rx�����Ӝk���ް�HQ�iD���C�[ت	�v-Kx	���/XNHt����6�&�;�>@��\{"KF|��$�~w���Ic[N�S1��w)Ė���,�<P2���t����-��p�2z��5J���s%7���=�|;i�'�����Q֋�Ǵ���
k���%�JޯU����Kw�en�
��J��'V�P߸���"Iݺ�Ζ�Z�D�:\}c�v2�A���jLӨ�� �k<���]G�u^��̔� �H��D-��Z�#�����eW����s(�pc�:s�"��N�*$�d��%h<��$a-^3�H�ܑ)�H�����	P��I�(T~~a�=���4�.W�
e�Lƥ�l����զ������Aƴ�*"|=CB��ެgv`� �P2��9�V�a\A��`�e��>�l�  v��G[W�YTwd�����o�DA{K��4d�����$�x���{]��8�W�.�ΟQ�܄1J��]�z, �֘�W��Ch#�ru5@��4$�����/w]/7-!����r�N�ر�;��w~��a�c��.p(�v�T��v�PF�fpޱ�o5D����S���Ȫ_z*'Պ�Xԟ[��u���ٸ���j�ϾC�� y�q<������׷�0Ly�zp�c��HIcWm62W�{��������� H !��O1�Ѷ��"O7|�B.�I~���n��""i,�3щ�ɺ�{OtN4?��2U��?"f������1[2�F/ʪ�q���ʕ#�CuPT!c׸���d�e�Sww�;��TIq�2�#k��K*$����PI���L<��3#�}�9pz�GM,�fww�?�E'r}�'�U㽑B�G�/	IR��u˛.�.̀Ḛ��i��X�Vh(K{��Vt���^[q|�q�O�)M�ATs��/�8�C*L����M�u3gg��O�����'�恦ٍJ;�=3���I��6(N�)��]� ��:U�QfK����J����qɮFDV����"�efܟ��$�0���6x�6�/��?=�`����S�"��?��w��yJV�i��ǆ�ŊŷX�2%k�n�)��f�:��&ХcU�siUrN�ö���:=��F	
J~|���l>��tM�5�����u.e AV��+�tږ�hx����(�X�ʙc�"��j��"%$O�y�$�R��El�E�KR���D�( ��wH��y���~�rg����w�on	�[�p���3�� ��ҳ�Dp�xz+��p\���!Y�?|�eT��A5���|�qy׋�{B!���PI���2P�8�Qw.$��h8$
���ZS�Al�z������:��i��I�5�K�b�F��ȴ��N�����<�d�&�<�TQ,[��^��p$��+��ń�ݿX������:t��"������.�9��e���0���<�wm��.n)�
�R���f��H�E�/O�ߥ�`p4�BP�H�L=F�ՒxJrj���
˵���w�u��F�Đ�:��2!H����ƾ�Ķ�]�x���$�V��`�[� �8@e�r
#�ʽy7�{�1�k9&�������j%I�"8��&&ԥ�������+#'x}V�n���_�������i��Q��QAZ��ݩ@$�-+�r�;\7���iQ$���b\�I����,7�ﶒU�0g������X�;HW��o.!(�#��Ô�ZIy��&����>%�&l�<�>����?	Q�JM��CY{z�tOY�����k9��G�f�=�/�E@�#Y�l�5w@?����6�[�#��<9��iHs�J��U��Al!,��"���OK��(�\ۇ�V�}��-��ǌb�ƪ�[��U�$�ԯvŨ�~q�L�a.�UJ���cD˲2�36�3�ƿy3κ�'����`
,Y�>��b.��R6 ���RiV��dl_r��,�]	Bb��c��cqy�W��4f��g)Z.B���4�oW~�3Sq� {�5��7(?�+��'�MJD3���#���d�LV��� {�qxՁ��5��F� kֽ�kRԜ�]�D�@.�=Ps0�CH���B� #gc�T��J��(�(s|� ����S\P��{�8�����n�D�LR�?����IU�JP����l��8a+�	!yY]C!_�����!S1��r�A�v'�[���~s�!�"���*���Ywt�<���^���v���1C���Q*7ho�l�4|�B�^@�OLaB��-{K;���C��;�A�LG��zz�e�X5{zQ���d�a��;�=!0��{��j/�Kp�y�w�7_��$?�s��(�幁��%Ҵ���D�!��6*�R��?-�SxY�oCD��ĉ���=�� _/¥p��]J�[E2垪��+�uږ�p� �Y�8 &�I����`�=�d��f�G��b�/w1�W��"|�_K�:3}�V�5�s@�Od��¦i�AG E��1,�@^�#��\��X�aIj����_5��Wq��P�x�H�s4k<��V���r�!�o����`��?٪�TU�J]5`.��	��UET߁��<Nٔ_w)؏��1�k����vckR6rt(V���H,�Z�}��ƕCU�a�Ո��%�4��;b��ej��
�E�h7�W��W� �����rvf�^ǒd �q�������w%9�VM���N��r>�(")Q���~G�Rc�����sŢm��}#Y�������5�<Q��9�X>��M�(�nA�y����Л�[Y-�9f@�6����DUɭ��q����R|J*����E�%�_��k�r)�Q����w�����)`ym,j�H�a-����2y��l�7Փ��P�)�z}�9��D!��l�|~�!A�ى�S��Oޤ��-Ҫ��l�>����4����zZ�����Ĵ��&SB1+�ũm�-e��.l���p^|S��E�4ֱÎ��T'�i�E�&*-��7���xR�^�NQ[O�U�0��耏��#�G.�h�f�����/��)�߬�5����S�_������]n8u��:K4W�2��ӸU��
R�rA�EO���#�(3޳�Α���L���?�!�2�"6�d/��'�,���KXp���ih��U�t��l�R�S�������0Z��6� 0iΩ�a���W������Cd$������4I1�gC�U�,()����C4ov���v���+��u�wO�]:���	7Y��xy����!�ѴZM������eV��! 6C���r�4!�q*��@�1��	mvtj+�S�eu,q�[eO�Oŧ���y�c��m���M�\n=��3z��c�݅/��L�MK�	ןA��~ѹ�+ Բ*k����E��|gt-���n�7	��
�9�͓+��y@O=*&e�W������`D�Zy�����7�`1���Q�]bC�--C.�r+� ת����U�ė��UG-�\=��y�C'�"�[��C(�$�2����"��T�v�/|{�;}Ԫ�@����w�!�k�����IL��5.p��m��*����u����T�<�E�L.@I���X�{��|�zg.��L�.�v���I2Y A��dt1�R���6Ov�3���0�h�a]�p9,zu6�{o�U����^zT���� Z(�=�X�(Q�Y�l�U�1�˱m���O�-�L�sմV�У�4Hc���G�1��՜eeS�P���%���q��Ty6s�O͢��c�
�7��O!O���Z��DkD�p]O>0E ��uH�l���BS5�"�r�7q;��{1���}���� �!����c�]�8C�^�]��%9��`�.W���;R�cx;
��}f҂����̸_ۙ ��)_a������dE�0o�{D嬡6P�!,���oeC�gx9o;�.%���f�q�J�W=mL&�{j�3�J�3���˯y0�l��ᷴ���������G1�GJT�Ej�XwN�d>ň�2����c���8��*m��sM���R�:3F;|���Ȕ���������4��雎9�j�7ܘT֥r�������g�t�Y��Gd�E䥍�9�k����r�}���f�g��V�t�c��G�y�<�̸�o`T�����0�9��n�ƸT!hh�cI��>���|7�(��o��Ӄ{�|�\8>�, �E�1-]���1�f	�Ǿ�6TPe�g�g8b�!�,M��mw�l��%C���R�4\'s��&6���P�Y�=����[!	f�7��m�\.�U騤�'�U����o=o�\y��T�u/��)��;�+�*��R��:��n��e�,G��s�Ďޘ�E=�������0�+�)Y�p�B� �\<{�} �S���B$�k1�$��ˀ�#h��j�[�{�H���v�ҵ���5���j{�L�ׇn���C��g�y�M�	�" �|v�RX��ϙ�J���.N%i��@����i��j�p|��N��)b��̅�=ڲ�o0�K�<�^�;g�oB�������FPI�j��F6�72�ϓcXk�P��js�{*Ðo��j��keu�T�\���yg�>�f5F�i..2SeS��n�����V����0ge�CmIt
2�w�XL�_��$ ��Y�t	7=E;�'��1��c��EN�Z2�8[���Qﯠ�$��+�B�y3�,R �^��9~M8��*���
h����(�2F�D�e�