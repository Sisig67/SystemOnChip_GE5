��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����P�^�Mqap)%t�?�&�Z�K�*���~O��in�ÇZ2���RG����R����k:�H����`�E�m��C�H��Ё�]]ѱO�UFH�Ꚑ�L
��"�0dF	�b5 �A��Q��+�	-�eD�4W!o�� �@G:�� ����Ͽ���˱z9-�n#��V�G~i�u^�L�������;�q�A�~��4�X�-�]Yl?/�Pa�����4ǱT|���G4'O;&�;�o�u���i~t��n���4-BǇ�aM�ݍa�ڗ_�bF�5�����
�s�c�<���w����\�_UN�΀'�D���+�qS�e-����@�\�By@÷�:K���F��W��MV�p'^���w}�#��
�VﱫIT����tL'c�>�F���b`(6$T�j�{���x>!���4f�R�;�'~>P�V���^�-x�v�:F�4�>I���Qn�0-68�jfb,:$�9>�X�y��?��vLr}p$?�Vw Q`h1���M;�qD� 8���L�-���1�#���Г#���J���G��Ș���H�������I7EY'��'ϝ1�UREcB鲱��|"8<T#���-dݣ%�*� �y����\��|�;��郫#������rC����n�D�x0#�z�wO�������F��{����u�$I8�m��y8�A�s���D�aehq�fۨ`.�
���zL|��˪o�I(��n�ZF�0��1����<Qdk����/�n^�������u�ڎ��$�=�[�[���F ��������zw KO8�>���X����$��]�JȀ�(Dm�{�̞1�ĩ���9��Is�;�)���D�˒%p�8�@5����,3$Hء��uEw5Es,O���s<�})�-��Y)9EW@��g����=���K<�)�k}A
�����r�1�c}�;M� Y��:�x!~��X.q�A⿓���R|�(o��bS�N�����$�6�-��D�J^KC��Q��A/�%��B�c��b�ϟ��Z���"z>B����wl���\>r�����Z8r�\��*��5���q%�'"쯽Kxid@�|`�\�5�&'�R�ѝ�1
�����-dLz�K�Мl&d���V6����X�sH�XO�nH�Ⱥ��r��g�2	�L��Icu���9�ލnv�N\�6]�w�+"c2���h�8F��Gƿ�]wR<\��_tnOI.�מ��|��s��4)p����������v-t�.�4N!�-��eZ�(�1��yv�~�㑹��Rݖ¤�1�@9��׸{A�b03LO�?c��\ ����]��ɶ��|2:�"~rE>!����<zoW��ؙ���G�]��}&�į\|����Z���K_U�_f׾�LȠ��
�"����p
�y���~=���?�P�V��i����è���sĝ֦9h`4yoJ�\T��*1k���)gW����3 XJb!�bC��j�����;L�SD[d��7�6���#�a�qMp���75�aȷ,]G�^��Yq��Y҆'�g�E�I���/���L����/��}� ���K��b}�b����؋�j���[8v���IX\������U�Y�7�#��+K-�tT.E�w휃�ɲ�~ARS٠?͉�T����b�y�XS�/? C�	�W���Z�5������!�g�K.h�&�.� ���n{�K������/
�//��w��?���jr��`m+�o�e6�ش�K�E���0��ˀl�}
����O�`Z�o2R�_�s�2�6�t�2�ퟮ�$xԳ�+�{Wr�L`L���u7�nr���J͑�H�UT��Ogے�¨�|.ekT��ޞ�^b�.�<'�������/�5W�!�u�4�9�\U��Ma>��đ�j��%%Z��Q�L[��f����֑@I3S���t�<.�/�`��
}�{�:��-uP��T.{�F�p�	W=8��Z�x�9����\�C�WI+�����|�\ɥ��^�i��%�Q�A0�2�)����}oa3`1o�(߄;^���=�g��99����	?&�w�[r?�'w9��@���(��J;�3�M��+W����w��7g��X�%��úh�1�P����jOt{q����M�Qavd�����zq�19DN�J�t ���L3^�o�L
s��V�Z�ƛ�6e�Xț5z;���P����/�U�v�w��A���|�պ����u�D�`�zp�����i� M�!j	{�����G�O9����0�OEI����1��}��DÐ��-�f)�:i<?h�T�n.�{� "gSԾ��C���@1����8��5f�����X{�z�bb�H&�	Ƿ�cM Ԋ%;����u:������fg���N������3�����f���Gt�E�i�csf�rnkP�y���T';���,����D+�.����B�;�FoxO�F=�s�X�`z�l,��iRѳ�G��"����C)�q���K>u�V�]29{�?E��8Hؤ�Q��O�>��}�!�ky�^~��.%E�ZAb$���\�Zp��"%̖C�{9{ *��*���S<�h��=����+n�N�Q��M4��-7�Huc�&��*0y��vؿ��W���o���w���l��� x�Y��6�@�ª��Ҽ\�#rsX;�:I�Bcx��S-L���8ؿ���78!�݅���#�7�ѹ<]�(��UI�Ǎ��<b���]VXt���,7l�^}���������y����u�ɹ��$S�dR��X�H�fz;L(3����f���$��\�9���;Y�v���J	6ƍ@p�|�)/+삤'��OV���z�i�Sq�\k�pѓ;&:KL#H/�rƷ�����ƛq��n}9U�s��7�MDD�.�}�+�r�$2˒1bSډ�_�WVd#�_����[uy}�pE�d�as�w�\�c����nx�=5mfڄ�p}Bq���s�����'/��)qdJ���d�*������5
^�`K/b��iRU�R��>��5�uiu���z����O����Ŗ���UM�Ȥ��'�g����"�R�K��>Tw�vr�w�Ϭ��U��˝��an֙�����D��'�5%�G}��ݒ��O<@tfrUh�YO��� �W�g|e�zqWw�Ҵ��r
댚_5�Ɖ`���*>��HP�z�d��}��H���S���� A�1D�0:p?q!�yֆő�\/W��s���a�!���m���l���^o �����t��[�����5�ՂE��L����k���o�o��EPe$.u
|n�$�2_@J��2��Ԩ>�Ǖ���(9Q�~9q�0l�{�f��O�xP��n�`�N�-c?X�8Q�j�,�.�߄J[�EFV�[f��O��gu���)ͽ�n��KT���7d�l�HV�aH�8���1oHe�wQ��W��o5r)ć�����mSd�����Ui��;����*ίf������c����d�iU��]v���S��L!�3��[@����'����<2���b�ʃ�6���N0��T��O?D��i���@54 ��M@�_�#�!!V*�Q؅n��A�	3�����N��1v@�P�;7���>/c󩀈*�`Ҩ�yک�����Χȣ|$(J?���ĳ��LF�����w�9'��bGV�6�iNDw�����4Mns�&뛕��=�$�{h�.��3 O�������
�g�a<5+�W�0�����7b|�)�jVX�5�_N7��1�Rr������%;Y\�BE�?���#'։�� /ٳJ�S-����e��h�����A h�B'�����B�Nu�Qިm��f
��$��|$*�	�|��i3-��C7%���W�3��̿�U<e�Z�Vo^�3�hPং^�\?�O���_D�EB���М،�_���մ�e�<�6�'���"bc3���A�]5\2�[.1r���p��l��\Zk�s���P�6��9)�t6n��'���o�QQ��Eҩ>㼽��[ .��W�%��؆J,�fs����m�Չ@����p���k�������e�/��t3Ye�/uƨ�Ѭ٬hŚ��&b�#����p.�̤c��O.�L�`�i���iM{��Ó��6�"?��Ķ2y�ԙ��u.�{�^���}�f���C��ػH�ч��t8;�'��rU���}V� ئ�KBI�iF`�%Fџ@{`���H�<��Ⱥ�2�C�<�2������t��O_����0"*�m�C�(�&JܘX�5�/������e�mM4�	7�b���8�&W,�O��׈�)%�
�bʎ����FS�K~\��Srn("K�NP�e3�g���'���
�<w��#ƾ�-F�u)~�vt��X�]0�9W�k�r�u5�}=5��?���s4�8�
�����w=�el�#j4:H��<I�)���a&{�e]���m�Hm��`�Z���l���G%I(�7"�������2�2+���������/w�)_�І�!|�4K�)1Z|�rY;7C����G���v�"MB6��eIW��y��k�i"�T���Ff��/M�R�
i�}'>I�u�O��y��ɺ���	+��tn�$�cM�}G��KnI���YKt��������.�XE0���=k����u&n�Z�r[���O�.��s��q�KL�ג˲�r"Ê	��Y2�?����lxvIq4x)oD=����i&�v9�U*��Rq�~q��B��?'�n������NN�<�A}���@0:GҐmg�-G��N�k������5g*�ӭ��K���6.��������E��nT.y�9ȴJ�<�@b��E���~�;������'�)0���˦��]ks Ʒ>Pӽ�$�%t��zn���w��9+�� ��� �3iO3���J/n�lY���14'Y���i_���ؐi�Q�$1rVoT���|c����,�!X�dkV���Iy�&��-'"�˂Pw�~o���|�?�U�G��m)x�
J�ʥq�]�N��-�gˮ�|G\
{�{u��߀z>c�&��҅���Yr�a0�Pe�R�o i��}([c����� a	�:y6E��;F{],�<���q�(|.W(E\(��hNK�-c	�����#r1���%ɥf+}�5T:��@F�2��zn�R�b��ui����⚬