��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj�o�v{'����D�Z#p9'�@�,�}*��[���� �,I�Q90%�ŌJ���_�~�E֥W^�	��� �njܰ/4�b�;��u>�y4���t�:�Ua���̹�4�D��jiņ���F� ���5'����*ִ+�?��Z��tfI~�M�{:�a�9N�o�|^[�XeV⹦����B��	?���^��.�	�i��Z���19���QS!�H�ʴ��#ql�R�΄e�t��uF�� �s���e����h�t��?�I�Q(����%]{�TRɤI�0�&����26��D*rVdU��1`��f��rj�N�0+�2���V���ԁ�)��Ǆ8�ã��'R�^�h��BX����`7&B����
�^�v�^��W��m.�����o����c��X>�jhSy��K�i��v�,\�-�|�7t�6����Age_���M�n'��U++��c��_9����8�����Y_�G	hg�`\7�c���G�����Ȇz+Tz��B� �	l�7LX!������A=��'�V�ɛl)Z̀v��ّ>ޯ���&��@)����H����.��gy:x���l� �?�^�D;���d�o�j$6��O�Bұtۖ�d*s��כ2���FUC�V��S(x]V�Qγ��8�	�>je�vL�=�5��/��a%��LҰf���	꧕Y�O.�h��୥���<<�4����B�/&�f�G���֕N��'��M: � ��҇i� 0�[��� L0������gP��S�������FW���G���h`R�Է���n<l�J@�(~mA���v�.'�^#we���\X��d��P���EH(�]�]XsL'�/'ߣ��X��b����MGz
=>羂��㚣<�~��,H������{:�P���<2ל�(�XL���]��>���B(o�o^�!q�F,�v��7�