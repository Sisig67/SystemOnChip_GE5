��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj�o�v{'��4�4N�m@b{L��� �p]�%F�  ��q��1J�F,cjjffa����JK�a<Lw����!�!��U4�b���������7hJ4�c�.��,��$�]��oR4wǅ8�`/{o"L�D6&��]B��1�����T�xZ��"�GS#��������<(�w���鳈�������GQ!X�R����Ԡ�6�����b9*�l�uJ=��mD��̞����!���iN��#x@a��fG�_Zu����Vcb�_��]��{2�-����!���HڄѰ#��x`CC/��IF`Ycyk�I�G����&�B|��^�e�ء�p�0�΢���s�֠���M7��c������(m���j��Ic�ws�Xm�q�e�C��΁����|���Ø������∼�n��ư$�Lq�3 �����Y�/����ֿnї"�i5������Nx����F�-�U(J��ݚ������2�VV�w���A��N��+
S�w������rC�^�5�[��J�!.�~D�V!�cf� -@U��
����)�g�@��N�>yR	�&��]50�� �W6��_�r��A����F7�7y�n�
"� cz����cN��{�:I- v�y�Ͷi�~ŹӰ��6b�������w�!���*�6GO
݃v �E;ceL�iӁug�B�$����(�k����FF �9���l|J~>�W9L�~�.:��:�$X�
�2+�k��k\��"݆�z���2� .�.���h%^���F)��#��xuV43�[	�v�y��޹�#R��U��8�Ϯ�;�Z6�d�_�q����Ǹ>�χ-��nAIǌi��� -���G����U�d�5H�<�6�h0��*����k~��9P�$�`b��b8�~�l�:��Ů��,������a�K��+ؾ�\ �޺'o�l����-���Q�Q���q����+�I��d�C!�X����5J�M"�;���@��-!$R�0m+��%�OԒ�6e��c�
��J\��yN��5��o� �9n�1���յ*�Q���zP:��i�¤� *|��HWB};�<���eR=}h�]��E\6.�Վ�3��!������l�ͅ�0F��I���Z��n����*��9��T��=��lW�����1��l�m
O|�VBM�
��	O.t{�C�I�}MXr���Tn��w�#�?��y�)z/���{X����vI�Z�������Du����V:N����Ӄ^�-Iu�d_lh���`G�V���;�z�k�U���t�	,��s��E���"�f�ۖ�|'}?�L�!��+���0T�H��v40%�i��Q�����td�܉��W�,�����P?gK�|tR��6���K�rb��u���>ud�<Q�|l�( R�[@.�ަw�ս�����Zj��]l3�4n�眿�Z�A�.���@Y}o����^�D�K�3��� K�u����O[��ư��+�,\w�nU㞯�{�������{��*+�P�S��������`�2�5�����3B܂P�x3��pJ,����e���N�z�0P�����i'����TYcg �a\�OZ���x�X-�C���rַl��eL��`B��C7gLt�Y���`�G:"�e�R����l���V�f�+�8,�E.�ٔ�
�l� ����8��'��H�(�Ͼ�/Z��CaA���ΡCw�
�SUsAn�"\Y��&�ƞ����}|��=�D!�oG�I$E��R�3[Vs��la�N\|�D�TLM�`"s���zό��5[yxcF� �?jl��֝^2��sqxy"	U�N"9-N����˃�B� kл��#WUq��z`ة9��Q�ۢG�g �ߛK���&������@f�`d�5�tSgz��J����b�������[�&�=����������H"�v��{WHUΜ?:Ϭ��A��n���J�K�2���3c��5.@�	�^f�W u�	���ՠ/���N�]FִJ�9��A؀�z����	q�ę!wF���4D;3a]�KnՌ.bfC�;�v�QhKaq-���V��{k�ăo.Ң�G1:I q�A&n�<b�F�G��e�O���
��1I)�/c�z��H;��`-tחxI1q/�GD�~�|0��E�j�����ϒ!���a6�W�nJG��Hd�X^���C;|o.\�Or�G鿀�����z����˽�F�T�EE-1`����(�@
f-@?�mb@�J}jW솔SaUB��!e�M!�d�(4oS$%�RE���Q$J'�ļ�/jۨs~?�a��)�H��m�i��gv
u��`����+3��vZ��=$�ז/iH� �~�̭��B��Q�^����!�f�f)�b([�fS���8��g����GR`'�W�<,�鲻�r��:M���_3͌\%�����3v���1L�2$ffA~�`O�v��I�%_f���i`�y��S��YӺYV<_�ʗ;,FJg��St�3�wӘ�p[��o��t��¡O�z�8��v���xF #��Ԙ��*hD�XS�+2f �Q�!Az�b�Qx N�F�`2m�>��٢����C�����ƶ�`{{����D�z>�(��(�R�O�?��ӽ+������3z'.��O����+Ԭ��J|��G����o��`�q{sz7�����Kc1]�n�cȉ!�<�1��58��w;:T#Ɔ^�����N�
h���)��V{Fq��-^�_E��M�-Xئ�oR�f�A *���$�����y򯄸E�=���HCY^%W�nv��-R��MSR��>=�r�v������-f�;7�������9��2�ӑ���w���r���:t�C��i�6�m��SbX��������t��9z�{�B�p���L����++82O�+7���WQ��-�,�3/�������D��#۽`�!�?$oF�I�vΛ���S�I'�3v�)j�,��>�{��ޡ��U�?�=D�I�L�=[�O7a��� �ıW���2��mG�� ��<�a*b���)����$�w��=����Z��<�C��Tl�G�eʾ�޵N�����i��1r=3L�*q���1��؆��Z���J2�\�B*�E8D�X�D�P
$�\�G 8���(�$o��4�O�+M=e�L��JDy�*ZDWZ��x�kIk��J.���e��0���߸ݞ�V�V��o0�����|OFцvӢJ<rp��dj�.s��ܹσ����~����%�Y��A��$
>��O���=��XB<H���M�W��$*����y�Z�9���W���'����S����{�H��h����s�5?��0��d�c��71�\�ڱxQqe�<������
�"0}�$�7[�����A��b���y����9�ы�v�J��1vI]�ye��o��0E��!CL�46\{`�K�j�MH�zq;�y=A4��b��<�o���k(}�k��xqp���<l�zb|�"����h�i��;B�{:�I,����{�;Ŀ����:��Ӏz�l�����pU��7P��@��Q9�A����,��C��Ey .�0�GZ�,	�f1��O��F�V_�q�Xģ�����_}2R]ڟ̞*]��� ��wa�[�L���}�z�F
1���n"���՟���Saǅ�6�`���:)�r�z�:7^etߋ�`���q�XЪɲ��aw/^��+Q�<���Ut�p:�I�4#�N�%1x#_�����9� ���翐���-)w�9GQ��⾝K
 ٌ����ܡ�u�Ɵ�{8"6	]�X9Q	؇��I�����h!��5/4j����Fp�:V�\�I+y���&g��s'�fp�+�T���L���Rn�>q�GfY +<����ي��zz�h��jjS��� �=�G�|H6R�H�2���O3q_׌�-��~0="�%���J��(0�^Nģ��߬a���������`���]%��a�k�k5 �C��ӂG�
B�<!9YJh����Cf�xΎ����p�O�q�n��(h-	�b��Rэ��MY����s|<� ��P�d���i�陛P�=a��s���v�O��t�,,o�
�е�@-��=��Y%p7��{F!�0徐H�Վa:λƁ�lk[���K]�++,��KɜD4P�0@^�z��G.�,y�["n���\1�5��@g�O@m�F� v��c���$Q̀�7<�i�gR=����t)�����5G7��{�`�n�w��l�/�0�2�~�NƯ) ks{`!� h�+x:��܇w�Q��ee#\�6ꖣ�'��(��䰱�D���	i�Ο�ũ�