��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���!<So���2��E�!�7���feI�R�34�F�\1uR�XO.P㤳��"����(W�����Y�us�'�V6g{���/�Y�^( ���Ne�[�����8�1��{SZ�k�eZɇ�FUHn�i!�kO����r�o�40e�@�̺Na|�g|�O̲s����_�oW�h+c�	��x�1C5�]�`��P�#�Ι��;<��C������^c�4�\us	���S���x�~T-���]D�lK�c/[G(+ف���j�H�3!`��|�V�k�)j���Rrj������+!�m�iS�\�,�D nP>�:V0�(�9��O�Y����m���7Ӧ�J�Ā7��-�o�6���d��iP�2I��5����^��1֐쬳پLƑB?�(�x����wj�j[p��ب�Q��8�)���b' �{b����Z�مIt<8�3�\;++�Ҭ���7���$5�?��Hf���*"��6u�Ea1�Q�g=�f	����%'(�l6���g�L�YG9�:x}�� ?d,2+5���1;T��U��Kڐ՛vN��~ō능���d�>��$�s�D�Kb��{��V�L����+��6pM�ld���v�0f3���w�ہ�V����W��� TB�Ov�4T��9k�m����Ҟ[Cṕ�Q,:/I�ff7M�d�$#*�=չ/Ȋ?@O����-�+�g`��0�E�΢f�Ր�#��l9LBi�-�.�{��޼W��������Jx�a�8T�r���ŲG��@�.�f!`¾F��^~�G|�v �FLN�j#!Mʤi��ɘ��R�������L�"��[�V:�(V�R�Н7�i&O��Q3��������>ac-k�cq�"B3Вa���-D��+�;�IYd�xޱ�T��F�A��Ji	���π�[�>pE�����ðh7�A�P5�f7������:��_m��\󔊁��?<���5|���b�P$1u� �,�U�����Q�	$��/s�QC��Tb�����nO���n�E.�|�@��}�"�^_"~B��F͵�U
�Zյ'��^L18ik?p�:�yo�K���&Q�V��b�՞�	�Ja�2��ň3�����c�R����k�����a +�M����,Y^����>b�D���Ͳ�J難��e�;FH���DA�ΘZ�K�\a��������w�u�ʄ�9^�H�Qf]GZ6�MI�"�N��	��, �����u`���L�[��UG+��a�HE@y�L�eM\z�`p����iF��`o�A=P���r8����Ԓ�K&W/�O�1�Y���[V�<y<Y^�±�3S�e�����j֬�\ML*������3���}�	���+L<
��8�iH�Ɏ̇/j2��N)��\5���gS�x72,q�/��Rw�9׀s�!���8��rt_Β�H��r
:�J��z�?�I ;��@�f��DTv��>M!�mHPDR
���ˏTC�o;Yo�%o��X��|h	����Jqx*�瀗��c�\�|�c̍r�`������:��;��b����� �=�+7�!K���[l�A�i�;�MN��J�/BX"��NBli-�o� ����t�G��T�0����Ej�s��E9Q�y��X�N���|��K;�t���+�xnҡ���{�a�.ue�:A���&�U���g�1�����;XBHn$��7T��2k�4�WI�*�B�N�>w�iP�-�=.� �`?Q���?�tS� 9�j9����Ӥ�9!�D��}�au�b��1���UD���O��	̡�򃵏�z耗���K����d�d΃�q4#��;�<yEy�0��-���%Y�#����D$��ӡ-y���Q������Br'��$?ۂ��N�q�eD�� �,=k�g]�*���<�E��Iy	��� (@�a�-�����:�̉U �s94���|y�"�J`� O���B^��*Z�uD]�_�Ÿ\#���v`]�slЀ_�~"kՍ���x.X � ��@ ͐�t�z��-4��`��8�X0���ո-�r{d��>(Z�>sVp��՛�i;I���2�m����,d�*{N:G���8��-�ٷ^�\�\�lp6	{���e�Ag��G	��:���,�7���D�o#���؇�Zo����G�޶Ym�;e���{&�^ H���)��I�ϫn��A�s�&�
�<�JS��������M���m}���!�����Y_���Ը��wI����Gha�AJx�_*����R���@����ke2�3v�.į�JȒ��������B�Yy�~�,�����[�����l٨Z�:����=����}�wG�����CN�����-�Ϧ�ȵ������f
��5��]��1(ǝ�B�����(l��N��䆏+L�[Jp]/Ĺ B�J��s4K�����i��N�S1I��+i%c�(��,O�!�!��
���s�n��8$���Ym� �R���fy#\�qBd~���8-���=m��A�� w��Đ�4z����-bjٸb�&�gp*���Y�� �����>j�_
�u�t5��-+��Դ��tg?dB��!_B ��B5Z��u�4V��K����z�F��L���~ր��������c��/5�L��1dŘ	[�(�3�7�
K��+E<�8�;�D�`9:��HfO�j]��U�'���ڪ4�_SM�Wg�2E��Y{���"l������P�$�d!��p
!��&w��ȸ��j���}h�k� ��4M�T8�l�hLPQL�d��Ǜ|{I;�=3�LX����2�X�R�e�I'K�l�������ۧA�Ð�R<�m}�m;�J<nE�F-��	��K�8���X`�N�ϛ�80�֥3�f�\�@|����21���n�2(K�é����[���������7�,p����8�qݠX�"Mi��G%���x��9�1u�~ǡ�����"���D�� TR�L�~�|n4T�ӟ�jW�0E��T�֠^�C�v�)���P��F���u����9�#@�V�;jq^F�m� 
�R3U���g�D��� Ե���Q�& �#/C�>���tz��T��q�/Nm�g�\�+@y�;s�o ��Q�AN�F�^h�nt~���Yn	����N��Ҥ{M]:6����V'wj'��q&^Hlv�,h�R�6���:"�3V�^䋗,�����/��ɛ`=јj�h.�la2�W�{����*����F�.�ӛ�B�Z���EP�a��2!,K�T9Pq��|��3/ 3�E/��<Uɝ�~v\�m��ޛ��J嫯Iٱ�v�r�[�*Gb��|�%�.�C�;��~W� r4���� ���Xpd!��v*C���~�������
`��IF�ƻ3�!��4ė��3��P�b�W��ƫ���[/�*�F�/�����M�׈�\�_��i��z���^Q�aE��$I�K�U\��-Oc�KJuͶ$,2Ōl�44���a'�R��s�~>�p�J%ڴ��>�Z�AЂ�H���<jP^uj�ybz��"o�	�7u��̧��Z_*w���Ihn�q{�x��{�����6��L��H��+���'Ě?���JQ�}�;�w�L��JS���DV�t�K>�ڡ�բW@��ɗF��+(?�C���t�G��ߞD �:�>^��𣷄���Q�q�T�=�~�m�`�#�ٲ@Ԓ[8~�i���xOOL,�A_�H"��E�J�$
n��t}zP0/l�&���ic)�ƞ�
��hx�n���Ň4���=���%�,c	M`u�ޗ��w���j��{}+���m��.��f�eǐ�m�,�3��W8�/�V���N˥�/��ͻ�+�^U������g#J	�U�ٓ`�`����&S���D�|�LJ�+�	�HN���D�=O����1��X����7IUl Q%Z�t�G;��D���8�����%G����	�|���gb �2�4ӎvoOb� _ �Sp�6PeC^���,Ǯ����x�i%�Qw�R,��l5�P}�����a���Hp�s� 0�s�3��^����sdZ��Jp��e�0y��ŷeȚ�������\���}���愐��?`�r��� \-�����hԣ���8�_e4c�vu������G���֡�J\5�E�7K�/�����d��C`c�u/_!5�*,�.N �]=*[OoQ����~suw��ȃ�$����hWF��U��T��?Ԃ>�~i��:�j'�%k̉���ͣ�����i
�nD��<*��}f������q���F����vD���ŔϼE��6�9ji0��r,�N��O�P�K`�.���4vn��[;��r�R-��+�f�_�LIe �~���tB�X#�g�}�K���� Ss1c�\����9S�.����W5���#cs�D-��/�.&�,�7�_�����TH�=H<��s�g���Ѭ���ޏxx��72�9��[�7�zS�N�mhP��n�M�;���z8��K�>�1������y�]`q� o�axgMu�V*K�8w��i۴�4�s�����>$3u��Jݕ���Z/*�x�3�A~؍
V�Oי�qO���D�H,1<۸�+�T#|(���l(����'O��q�hFN��+�J�C�<�C{~s�h��1��<t�t�`� B��!۸�4�2����ε�tM����Y��
�5h�ydNm_�s!,>���2JQ�?0����(�%r�9{�=?p��ӌ|�����>!���^�g�^q��\	x��S�"���F�q��`#�C���̄�'#�Λ��dK��>��C�������h�D}mrot$�e]BW��'��U�u �b�%q=F;�کS{�h�A}*�75��w5a�&k�$�W�����ٙi�d�waN�:4 ��J1a���<P��F�0��ru�O6�0��@`d^�2�R�)27Ӌ{��J(���`�)L�}��֖XC�`w�A���v�Ӗ\H����0���9MhΎk~�ry��[���|�u&�Qd�,���y���E��;n/R/̢���0��C���1��\��ة�����L�^LU�9h͋|�.���:He5��������V�ȑ��fbC	����9�.�H�ԉ������'4��VקL�m���>�M8/lV#)GZ��#�̳C4�B����A.�Z���}׏@����w���|��~�a���֥#"o-����T �V�(q5F�}l��x��?�!Yh��f��<t�d'��C���G`�m!"�Җ��yMs��}�Ͽ���4rߣ�!4_���%"��bR������
[ʁY�9���`���}K� �ǲO\.�׹���Ft�y�!��4�K�J�??L8��]X&6H���T���?���&Jm�jGf~���+x��g4�C�9k6�l�{w�y~M�a��Y����bB<K3#qnDϣ�8�T$XԼL@s�6�}g��Ҍ����&IGؔ��gЌw��ѯ�S8��c7K�ع����l�/4�W�eSp�
6�f!���3+�!��8��{�5�3h��L(�YFH�fz�2��^��A��ĝ�2�i5�d�+�1�̃�h�h�5��@�))}IQ����unqLZڟ(8@�9.�/��l���;��l�lo��`�RBc!���w�Oo�sN�3����0;_��s���G��WH�}?).�j�4���h+��K#����������fT��)���hLl��9�T׮��7v�^�D�t����u蠊 D�*�0~;�{���%/)%�b�q�D\�X$e����!�&Jn�g����t�0���VF�	~�s�ka+1.�#}k�T�Q��Mt�i��HΩ'�Mh��CVf���P��yHݻ��bL~��!�ԕuyP�;H>�N�I�H�u�p���ګ��\=��  ���O���@3ʙ�kx���Ju����2���ɲS��3N6yS��X�ƒ�k�YC�t����4�!`��"�F�[�m�+�˟�	cW{z�V��(޾ףvzK>�6�Ȗ8&�4"7Y99���Y�r�sи��z���~���L�;Y�����>�
�x�`14��V)�"�{>2+�@W�xgS1��Z�4�mxo��π�z��Z��%Y:UR
og�gq@/R���C��Q��,GI2�®�Ǽ��R∓�&��z8�-��K��HP?���t��_��;\�D .]�_�򘌪`� B�9b�4OR�'��#
̀X�i��<l������?��.ݒ�I_�A,20��>	L�g_FO��D��$��E�-QӞ?��������c�1е�t�$i'07Y$�FS���q��$	�-�o�CM������F��8%�����UȞh�k+�t����
)M�5��Z�tD�����>�~|��"��oH�pI0��!���LH�zj6�G���8ZL�T)?U�O��*֦��A�V��<x�9.��sճ�9$�N�࠲ Q�OԪ5L.��=zb�է+���O�������L\�!�=3�߈H����:AK�CBX��2�y�{��%VT��4)��W	��M����@\���o~�Wy���r蹿�hmJc�vb�W.���ŲV�R4�
�喠7��)�U"��ޱ� �#�,����0*�o��+M�0R����9��O.A��-8��m0�v�Q�
h�M%���>|�2�����9cZ��j�<#�;�J߄��N�����ȩ��_��7{�Aڣ��a$�/�j����G�j��݉�R��J����
�z���
���#zѻe���_tJ�f���d��'+(G�8ݏXN8���Y�h��_��EQL�W��`�2��x䋛ɨ��*KL�U��&q�N�o�8�U��w���z�?��)�3�gu��n�s[�8�ˏ^�˺ �ה�$A����MMd��9Hi��%S&"�͋�f��7ˈ����Z��#L~�C��Ne;D����.?,JHk�צ�$��o(5�Snt6ec(^'|p	l�!�FBQ1����F��40�A{ߓ͛�0̝0u� �k��7���(�Υ�c�S��X2L�֮�fJ�-���Q�op6���uQ����L�]JKep>�%���8������y�@����<FVʼ�t`�.Kz�uP��?��WwQ:d�#�(��Iqtǌb��~����z��ԧ�AF>&�%�{M�]�N��"���C�9؁{5������E�T{����DϤ���
���sa8~�oS��CA@_��>.��G���:y����3��OdBAx��v��5S�J�E��R�@7ҨWD� �/	���!P���W�]2N^���G[?H��L؏|�/S���r��煣�50�:�n�5�K^�¸.�ci T�����s����-~H�����Bc�����.mJ��=/��b�ȅ1���ա�q�:Y��+��+O�A�/�hq��&Z!rs|�IV������k��F���$�%��X���p����ič�����r����R4��(�K�@l8����	)�W&k�S�G_��&���C�����
�~�ʱ��zl;��>}�޿�ft��qT�Ս��H� 4����u��?�aO�*7��k�Yf�q�R܎���1Ky%ѱ8=��f44�
�6�C�q���d]�2��k�t�`����o�h��L��|N)wB����ZF�Z�n�X���5�A˶�C�h�l�acr�q�š릇�����i������t�K|Y=�u9��*i�*7��`b��>����-�!q�p����Q5�({/����%�C�Ϊo��6�N/[!��U���8d��h�p�B�W�/��O�����H<�$�� (��hT����nd�'�!�%�������NA�t�_���+�'( �G�3Ĩ��<g�;b{�Ҕ�\�L�;�<8�a*�H�����=;���l�ـ:������?�����Z�M�I�fA3�6"�M�y�m�E����Mu2��X�$��Xc.��DUh��ܫ$��o���]hm(}���b�(E�t�|�z�i/m�h$���/ED�!�π�f2~��N2�z�P��ͺ5�
?��]�W��4�M��F;�ϸYX��N�3�Wy`ǃ��9`��$e�=]�l/������f,��d9�:3�k���81��c��Y�
�S���J|0�A>�.�>�(�����R�T���0Y�;�	s(�C�t���>��˸�Y�C�+W��b8B���N�ob���~�P�W掼�x%���6V�]��[�����M��@:�䣁Rڢ�a�~u\$ۭh,��4 w�}D�e��&��8�'ya:���^������*�V�l�&��KoA���W]� �Gz5�*x����:1�M���Tz/SKs�6r��6B5�Xr�HW�<j5���j]��CW���+���Ȕ��'� 51�+Pv�z�U�mļ]tl31��>i�v��!��;��(�:e3X�������!s]��)Ջ�Q�E[��}�Ĝw-���$�	]	�w��*���~���k��s���fO�q{��/�N���%nO�7�yW/7_O��(������&��A=����.�&�2�^��	�..��h�����du�Tb���%��7Oƥ�j���~�ۚ�.��W��_��Z�߱�Y�&1�����2�`�����6�}:M�t�F�g��_9�˙���9*�{�N>�y�c#��y$m�3b��2�$��<8=y�F�^�֔�І��BM"j��4g�lX�S�:�P�����2>Z�q�f��|B��-�����K��޺_��	�Gݽ�`!�a.���ޚ����ܸӆ,�@Je'�������,[^�D���/���Ȭǘ�*�0�R���F�م�6�s�v��J`4��V��-v�5Z�Qu&�j��rb0y�=��(K,/��J������g����S52�h�7���ٞB͏�oxOaFZ���u �OҊ���D"��e�I#��㉠��/:�`�S��`L���J��5tU�l!i��29���71Q�����'��*��V�Ő���qZ×�ͽ,�]\6U���ui%�N�[D�_+"|��r��?
!Gp,�"I�QJ��y\
�m��2fV-���;��HO��~W����M�M��}��	7���Oa��� f��q)�E)��H����r	�h������x�3�i?�B�%�� O������ÆD�z���SS��ϭD�����.�r_Ԩ�U���L��	{�?{+z�!��乮��~��)CQV+�wn����n̛Z+F���]:�2�D��ރ��E�\h�����&ue���]�1dߧcK��^���O[9��B}F-M ����8�J��M7(�Sq�Z�p�I�ǍH��e��c\n��_���u@����n���l�-�ӽ]��UkCg�OD�i������w��|��"��e/�'���9�F�y}ހ�E���]����Y�=�C{�Q9C���uc����D�ԩ�O�VJ(ĳb�	�3A ��j/ϊLN�*1'��ڇy����\o�����F��`�A��t��j���SJ�eb��A����9v�/
�"�B~��Īp��f~ބ�]���S���gSߡ�%�^�g��%�" �ゲ�#��:������y2Ad�����f6	�Xí:�B[M�K�bf}G��w���#H�������L�i�X��g�]�L��u2O���}ݺ�RbXޖ�
WU�����e�4��pV���s��-�:(�XB�ǾR�n���׳��f��ғ��-?æ�+P���B|!y�)$�߀�T�Xft[�m����Y��Ğ���Tc�9H���pqI�du~�i�����{���HJ��Y N0[ ��@�-��`��-a^�#����?��e���`� ���3qV?
N�
3O�N8+4���P53`�����$��7|�����XJW���Q�;�C,j�j���僬��n�e\)�-������7ڰ /z4m:�l��Z�� Qm'Cf�~n������T̑�⪣��O��3���:UO��B�):I�3}�Ϩ�A�8U���仙ğG�P�\�u�9�s�J�dp����2�T�G��_�;qb����Ơ�j=H��N��:�BisO*���V �u8�'v`��7?ޫ�c��KB)b=�rF���3�P��"phK d���"����n?���pƣyb��s�x&���$# 2�:-]F��{�P�cX�ѽ7:�J8��1�?�¢s^��TʢP�ö^�Zc ��g�f��\�sI�W���3{i<��2Y�@u$oK��z4jxf�c�`��ȓ_%��D�*^��=֍5u'w���L�Y97B,݁���]]��Lty�j�Ĕȿ�?�#PP�|��l!��)5S������uō�N���]^���ǥ(�׆jp��-���KU�֫��sA���"(~,����0����-���B���e����f���O�a����R���a�G�Ng��H��3�>���k~���y��^t�3���Ց��Z�E������E��A'J�-����ps��'%1�� B'_�Y��cd	&�����Ӧ֞3?�vⳬ�����i�6�M6	S�"��u�G1�4�����$�/?��c�o�[��$�M�Z�c�Z�Hն4��Z�7�������,�	�d�v�����_|��T��R�T�m�Z?�}P�|I�}�!�υ쁋����9�����V�����ù��S r�8|9�*i	�M,"/�(����ai�B0N��j����� ��YM�J�wHB��'nW�i
o�jtj~���c7d���@J�/@���/ݼp}����g����P���I�ߓ�9�o�'��I?C��;���j���N��!Kc�7-9��Pj������ ��ƌ�'Vm��L_���'Q���!a*"���M���(�jPӹ�m4�7��|���[4��vb���ż�Q���r��$�r3��}�YH�S���:�����	�'wk~�?�ݲJY��A:~9�~/�7 BGɆ�6d�M?�a�"��Ѹ�b�����?�_�3@q
��s+JF��;�/���Sث,��G
��[��+l�E&?˦P�ȀGq	o7E�u��p1d���7E�Hmң�at�y�'}��X媛�+�%�]�PA��nBnt9������qV������V�9�	�6����Ð&�����w���m������Z�`��D��t�<��@�&�M����e1��L�)��ư�p�yC��ݎ�h���k�����j��4MO�l@�f��N>���"�-�V�FWp���.I8Vt��%���S�DFX?��~�|���:�5S���,Lgǿ�j�V�ufCpЭNM�T�t_�C����F���� t؁tB�|xΩ��j���W�sE�,(��r�G�V�R����cE���t\���X���%���u[#-�f�)��6Z�m�3�qP4��J����s�]`^Yɮ���.�9���6+m�UU���ȓ���t/w���Ӣ]�����,��sG[��[�[�s0�.s��ƝUs���_�sGx�B�&ϐ��M�^���v��b��i�ζM��Z߷؝�#,Im�Ժ�Qd(\G���4��'�5�M\�U�MW�g��*��(NU�<�<|��C�ܒL��eXD�e�e����ND�3lR�vѬ���MY;v��O�QT2�L����ߖ���)J�X�Įd�ym}��G"�:�#��*�xC�o�\m��=|ǉ���T/=2�y�~.z�:=V���^0���%҂Ɍ1XclǪ��M�n�:5�{!{D)AYU����FP{����#��2�?���HK�Ey�!�y�~�a�+�Wۑ�1�:|���b��i� T����PE�����h@����/�A��z��Կf8��*!z�=\���8������E�8���4�r(�O�ڛ�Y�������������,8�F��Q�K��O�n���Ka_�Nj��bv�QE�}�>D� ���z5��Dף��,�^-W|�Ο�&V_.�L�Cۋs<�=��cI+ޙ!��'��,�$ �p�.�Z,Hׯh�ܞ5`��b��]L�H��%�I8��FC������:��T�ʃ��<(3[�Cg&UuՒ�˻�;�����@��N/��i�E���XA5�Z�5ɦ�v�؉��E����m1��2hK2�d�����#�	���  �Ś�d o�'b�H:3_2�s��3{��s��aL�UO"�@��L&�z��DoE���]'t�����ڒ/�n� m��#�t'T��j1H"������ ���|PDY�K�t�����.�VyG��e�{o �@��~���(��Ԝ)وs� gLE�j��or���hS��e��+cl&R���-ο����W+�ڐ��7%��$|;�D�G��A�3کd���}�(�Wa��#"�z���z{�n��	v�v{1i��0�p$����V�?�d�/E�΀s�<��G�� Qg #gU���-`�Liu~�I|����=�����x��7�}j�3c�sQ�p��k���h�V�:z�`̿i����4���q��ţ�r)�$8{OaL��\03�s����| i7A��.�E�g`�μ˖������itu\H.��!�SJ����f��$�{���	T��yctR�b\(hcY�f�8��DfN4��H��hG�ps.��!<�-���~�y�������{��h�m�Aj,-��#^�Gde���\Y+����q��NB�jA*�u2z�~y�,��V����/7yz��K�Fis�����d~[�q�[ֶ!�ҧ�Z
so�"2^���ӏ��[��?��_���VaC2j�(���b�6W�Ζ� �`�Ī��I��L��~�ڰ/���Pe�נ�oy�o��QV�/�):���_i����8���g~����¡F6z�@s0���o�	�0ѐ�$�J(���=��ⵉл���UZA�Z��A��0� 5xc��7�Pl-�7�=)ѝ����H+�"����E�*�P]T�00��l��|��9�0�[ޗt�4�o��� ����d���`��F=�i:uL��c{ ���C.?'Mu8��8!!����r-s����F^8��|J��J��Oߎ���ER�5Er��h!��q���S���7���$���+(�p�}����N�#����X�9�Xl���f�ϵ{�@�}i�g������v3B��Z�{�G���~_��>���e��Qn]����f��>��Ӣ�f�]�i�Yh:?�c\d��B�+~��Ԑ8NԶV��k��}�CD��+j��,�"
��6B�.[n��;z��������x�K����M�uh8��ȴ�L	�F#i Te�dr��ok��F�	�'e�fO�0)���G_��K-���A��q������MB{RX;��E�s�z��u<�Z�k�8/ߡ��X�$�r�hH:� �������Z�t>�/Z�ꁖ�{a��1�ʻx����ra�o=h�Y��%�;`�&�wW�ܸl�+��c�� t*�a��o�[~�	�i]�q�8C�(2����|�>�_�-�6@����.�L���̂�&�(3d�([vW�Ye56�38�f��<O,�c���ߛ��� fbb�9�p��X�t���WL�G����X�T�Қ7�R��o����b��OQω��$�����آp��;H�f���3䞆�)�o2h:l))kR䞎��̖=��I��M9�>��`�
I��7����p��HT	"�]��]q�>��R4h݀����\��*`ɏ��s$b���gZRG���P�܏��t/
�5�9wR#�zd��H�ߐ�v��/�O(��L���@�@Ȃ��"4.=���-�-�6���Mb� ��4uc]+ 3��hm71�z�U4�?��TbK�;8��>Bz������7������\���F�dz��4�n�M��eM��5��Gҁ�%^$�9U��TN��� ř�m?���	e0��8Ʉ�a��w��A'��j�-t�8UoY�gJ��gc'��=��k������Cv:�	[Q�nZ�]L���F�c.ٯ��W�Aa�����&[a��B*5x"��3̛iE�ᗅ�"�1����,~w�K�];�ѷ�dR�p��� f�O���>�-H����\{5ͺ�������	����������HaD�t��,<Q�R'lT�/�C�mt���<��*�Ϋb�Qe�B�Y�<d0�b.���C����w���
��V ,n�!3�����3E�HK�cpw�z�@��� `��|���j�����"��a�Mq9�[/�?����^>q��"�]��.*a��F�I��@��s2�����0��ӛ-2y�������E�|�������R&��>���~��c�f���+UhHu�!ͩ�ÈEk���Tm����c�gл�f�ޝ������s�u���Z��`&�s�^�YE�~��m�g���v���
��*Q��u�n���M�$��e��Y��Ei��DYK{o��+BK�֋O�r:�:gć��+��D/���^d|:��O�m�Ugq��TyS	�k��F�c,yB�p����0�Yĺ�$�ܲN_E�󑘹��m�XM�����WP����B��S2�cvG�ke�
[���c��~��`�R	'��g2z����j�T��Nf1����%@Nߐ��e#��c>��Ntg��8���ߴ��è��� �׹Q��O)�Ͷs�����H���g�ִ�������!���cm�����'F�]6��0q�W�-{g4U���:uim�֩*����ø����6Ѻ5o�~�"޴�'�M�pev�DKDx�WH��V�n	�aV�Jh��3���suS����D� -�����!rD��/y"���ι[Ό���]	d�[Ĝp ���y����ȑtB��݈Xr�m|j4_���$s��2��ӂ7��ģӮ@��m6��ܡHs���X/9�·ځ��9�����֎��1�R��?^�������i���d
5��l���.�p�p�Z�w�/�K���/ڑ13���C>\A�v%� �˶M�R�;%e�5~�kΔ��(��e�(=fxY7G}"K���`ϓ�Z�+%WR	a�	�0�i"�V�ى��m������nLp�tH�|w�|9�B�)4�	���%e�Z��~ӣc��){��/|�e�HAV!�d^zM��^o�&��թ�r���/���[������}` (Pi���!�ٸ���7SK�p�,2�u�{�вJPI)��u���%� \C��^�1E�*9�H�ȥۙe����\�L^G��q�}")M�� :;i��~�U��l��/�`�󺔀�Y����PE$Y�7�	�0��c���i��Zؘ��vi\��T��%%L-�����M���8���"�3������{赕�J#��\�;X�l�V �:8Ja�M�}l~
$����X���y���=I��F�E��!���U7E���aр�r�@2���ɔd��Z�iȚT'O��UV�#��y�΁"�1�S�#i
_��:>�L�T�ȍ?�s�A��v�T�M�Ý���=2(���u�м��i��jU�m�����Z
�P����� ������~�%�͏��2�l��0���&���I�z@K�m_\i�L#f��/�6b؀��Ou�����	��x+y�����ͩg��b՞���r����t,{��t�>a};�)�����ES�-<��y-�H{�<�����.蚮_�u�J��hnpi�K��+�
�&��S
l�P��̅p'�r�P��^-TN�����!`H�\T���$Ԕ;y��18��e�fr�g���l�1�߂�v�\[�Ο	�4�-~��]p���X|��]��*M�ϑJ��`?��,�����*�#WN&*�����zV^����'��t9hl��㊝�_�?a�����_�� �4*�TOh}s=�_N���߀���c=Yh�?rS�q�l$� A��@r��pUC����/�7�toׂ�Ma�{��t��6P����/s�;�:�s�����ɲ�L�:Ο��w��t"�?o[�5�9� f&|��3n4�b7�����ؘ�'�C ���F����09_kp��Ki�� ���I~B� �40,�zG]\d��AмCa$&q��
Q�`����)՘�գ��7J�:Ĕ�>��K�,nw�-�x# 3���`샼��i�s�C�����:�� ]߁�L0��IE�X$I��т���ET�!>-��6}�9���1J��3ܰi�LzΞPT��;	���~���V�J;�XOM���b��

���꾬���??���a�G����<pj���Ƒ�����:<�h�k��"h����zK�6�'��.�5�(��'���V#*�ܡI��}1�h��w��S+ �v�'���
������u`K���������$�t0�����39eGҝ�
�xUT.nw̽�ٞ��-d�G�1ں�l`�5[1���S��PO5g�p���p# �ĩ��$s�������2�����68*i�#��ǚ���lr�P\�#����x�>Q�B��6�Ɓ�,�!�r+nA;�`��C����LO�ч*n>cG�W^�/�����+��a?)$��B^̧8��qL���s��C䤎֝ ��U�q5�b��K"�6vo�:jLo��uA�(p!�Y��5JNٷ~�Uj���GH]�@epx6��;DRW�$�0���HatF��0�{�q�ҳ�2��c1���Ĺ����`y2��oNJ�����4C#!�v1U!�l*�PD��'̔� k�K�"�����12�Ӯ�Fڑ*S?�\�9zO�2#Hl��W5�ܜp-�(y�#���J��\%��wl��ռ
}�᠔(@���A��#X��Z�\�30�uB�K�z�s��'��?.s ����W�i��UK�V��o&�N�B[¥,�@�Pb��pV>>̇�1���z�<1́�]�՜QY��QA����3��I��:@F��K��n�
�Pzw�T)�~V߽<D� I�َ%b2������ ��4�W���x��z��n�4��;���[6�,�V@��MW�.9;��,�b�sQF�͙�gLGR��o`h� 6:�$�qַ5&^a3퍘ھ������/*D�Yٜ��#&cQ���yhc�ԗP�z��$�^ma����A���*�̆xڀ�� ������Y�S�)Q{m���!�%r�M�A8�l �ڋ;����-ߊh�W����#������j����@�q�x2��.{Nق�e<
���"�AAaÑ��h�mI��!"� ��rH̼q)E'J�D�urY�N@��m�4ֺ�e�R�m͆˞� �̖���@��Ĩ�G1�Y��3� �����T�w==����c�f�=�D������cр(G���K;������
�,�+��"K�=�2[�
��(�q{��ti����!h��͹4m>����2�&�!�� J֤��K����:H��!0��{�{�S�T�O�T���i�t��j����#�Ή�k@���s���4�����Ƶ�Շ�)1 ��w�#}��p���xE�b�zȘ��A���U��+��{�QZ�q���� �u-%�j��y�����L�JW�m�-������ѝy�Ȉp�w����m+{��2z�8�����d��ʛ9e�Ufㅁ�*`l����@�4l�,:��AU��>s��syF�MN� ��nQ���j^%/�\���I�Cf�Ϻ?^��OM(�p��̱��`Fڷ����S�4o�t�L�f��f���t���X�l]�`��4��1��D��x��r��PmIj���/+"/}��cN��EDv�͐��'�3����]0G�CHV���6˦��Iz��r�	
���Щo�}����PF~��Ү�?2�m�Ѝ�e��l@LB8��i��E��Bx�=�U�B�b�9rh���̸�La�ʹP����w��į�=�Hc�q	��w��t�����҆����jϷ8�kziY�P9r�����E��f>���@[�Yk��x܃�G����oݘg���D�Dr�uJ�!}��CCN�����^vu��u�����]x�vp�~V�i��\x�Ww
��^�غ�$������6^�v��Q ��ؖ�������ih3y� �F���}�x��3��n��j��җ��#8�G	�:C�����o���NJ�C�8���01����M�%y	L�x��.)�~��EW�q�I�p u�L��ĥn%���f}F^>qHas��F5���QӅ�5ke�`��du�>��c1:@F����rڠ����t�e�D	�TRi��~!_G��s�o�8��O�ׅ^77�ѻ�aW
҉J��4��>��}���
gdC��'w9A����:�Ss��n�ϛ��8��3Z%_�'��с%^�2��~��\J�~��y�"�
:�j8;�]2��tBn�X��埖��g���Lh�#����.�����c�4��Ø:pc��Ί곰��x��+� {�D�cPP�MiJ|��k<n���c��uJ�G�^eƜ���T����q��[���#�΅��YǤ��ԫ�Fq�Hy3P�e@���5��Q'�z*�ɦ���У	_0�7�-�ԫ��94D#�Sv�&�ch(�� �R�0���1m�_�W�Ňё��Z�
���5W�eM#�j���vH(����5wJ�iË�NY��&�1�ʲL��������iZ,�m?�I_�n�����MC�ip0��l���=W�_���;��Im�oXԲO�������jdg�c�̨��v��%K�����B��t��k2�hcvN��9pUS~i��ɪ��E��P�������x�M� ��#�����1�M��)�N�A�9��u[�{�JL�?����n�$��Ǥ[#i�c/�vzn�l��8>���E۝����H��߲���zѰ"PP����Y�D"��'P���fw!�h�s���z���}`'���Z�N����!�xJ����h�����/�B�<�?���A~�SĹP��B��Vr/���5�)�e����_���J���<%@�q<<6e�_,^c������CS5AM��^~E�#�v�!kV�9�g��}��mc���-k;�AL�q����� ͮ��B.��b{���iЈ�:������X֊�J�4Ԥ��n�$�]��N�3�h.��8@j��J4Y�ͱq@c�8f�3��/�U��>�a����ȎM�p��3锓�CʝSa��K�H�%]w�~���taf������rh���5��0�����`�ߠ��^gf38L��')����
�5^ǭ�y"8���e��ݱ|�l*�Wk�������# �}Agp�Tzo�����ث��_kyY���[�';���^*�ǐHCB�#�l*RXTW�{�l�8dE�C��yyJk ]vKy_,AO��`� �"5
̶�iowChgujF�������f}9J�G�:QB9b�H����K��O�������Ɲ����FD�`��� �9X�"c�K̼��l}�k�s��
Ea���W��G�-�zE����M���4J[��� Ɲ�V��%�^au*HE�Ip���T� ܻIа�R��drs�%��M%���iQr�q/c?�*>���O���u.�r�[��1|��'��A��9����A2�p�ưZY�" �� ���z�N�](.���^�(���t'��G��_��Rv�&8%J�aA��;x�.�����8�b���rGc`[�~#e[��3��HijM�K�y�01��ly�{I.&J<��O�҆�S!����h�Y�}��I�	
r����#IL��q�i�c��+�֬��9c+�kS�J���i���Ċ4)�����A�����M	U �Z%�U�>�$�a\m���S&�P�ʧ;Du͍OG���0v���mc:F����L�Ɠ{zY�,���E+��gxt{X��9���gl�Ht�	�ȗ ˓m�����
���U����|��B��C2�֎1�#�YְN=(��ynS�L��/��5E+E�^	'�!�����Y95r�w�Xv����'`��^�]��-�`�q
P���Pa�%�|�/24�)+Ƭ�8�F���cl��F�����*B�/FO^b�#��ی.>��I��a���/ؾ�#��$d�P��ے��el&z5^9ق�B����Ba��.&h�
��go�Fq�o+��SD���j�c���Z�ɺ�A0�U7����W��]?X(}�Ν�OL4'�zi�Cϓ��L�H#)����V#��
��^!nH*g��
�X0g�cG%:�T,�K�P-*�^�ַ/n�g�tpK�ieڬ�
,4e�"Ez�����^¿6x�.�|�R{��~�u+�������l��5�l ����0�Ts0�O�|5�8�W��9����]z��B�w=�{DH �����V2�qi�r�:[q%��hyi���T9�_V�O���m�Z�q=� u�*dU8��lMݳ��&0'>⽸E8��Z�Z�b^o	�T��&a�y)KL§�I�c�y�������HP}��4>���D9���O�b�JK�{uf��$�v\ּ
�J΍\��6YN�kzs�)���_�V[�#�$��y6���mԁx��h����P������,�[)nI۫J�-��x��`�ܦh�L��=3ݲ�|�$�h!{{.�,a�s��c��:��º���\�Dw9�a��|���U�GeA�ȶJ�e�{K�N1��S�F�K���ݸQ9��W��'���WK.X_��m4�6g�����/9l}�Fq홵I~�6F�X��X�Y�#�Κ���:/��|=ӿP�9p��e:����2;���FV�@��T�
��1U�a�+3}�+	^��MN֊v-҃Դ�V�s6��8��W��N�v��۬�H�a�)H���4�ZḰ������Y���U��(���Ky׌Ѽx	 }0�-�!�W�g � V
�Uw����������4	��F���勺�Q��[<X�F>�X�/t���8�j$cqX	JF��2	��f������x���x0����Iv�w�	:��~�)������x:K���(��Y�~�i���v_��@u�RW��#y�9��l~���*���� � z.�q9љi�D���#࿷��q��֛�)���l-�.u���� ��ɔ@�X}g�nm��` ������."�k�M�����RP��ʘ>`��΁�O������<X�wM#� #B���bB��G*}�����l��R�ÈPj�{'�3�w�Iˤ�Ё�kQP�8�p�F���ݍ�Ao��Y�%M�[�WV�� +C��F���,������C{�u���m�K/Ƌ9Z�����8"�	i�{J@w�'�^!��*ugdr$���lB�Ｆ���{? ��������45�Ŧ�3��4������7Jy;�ܨ�3q��&U��"��1l�}83��+����V5ػ1�2�-�s}4��zH�	*X$�����镼x�&�]E�=��,���ٙ�V؛p@[ͱ�uW>7<���g$a�nl�6�����;�`$͵�CfԦ_�y ��(; l��3�Mp!N!�B��!fs�LL��=�n ����yݶ�HA����>���_�4���"��;V���'7��D�w ���)I@L����V��)����='�vnm�>CbNq,�U�#��ڲqYvMUBh�X_�h�Z���w��JjO��OP���O�:�Xf柍�4M���׈���^��~�v��]���2u0G8S^�к����?�ȼ�_u(^ ��>�v~�?�AE=�x�tT�W&�O�H ��dps��S�.7��]�/ޛjg�����=LG���[�A)ʆ~�p)� J�`��^A,F�4�س*%Q�J����3�B��Y�(�6�9����E���T�*��l��Q=y8	����F������a�cGoT#�rz5ѧ�L�9b;�NrlO;�����|���j*��<ϣ�6�X�������Η�̇��&�~�K��^���{�%�NL	S���x���>x�n���-삖�s���9P��Q	D��]��?b]˛$ ��H���q��[��[��(� %��AP*e�ck-ó�$�шI �ZV����g��L}����~�����Ђ�Ȝ����}1�oD�oohy��ʥ�3薃 �b@��-17�(K;@�@|}�I�����!;Ɋ�pat���f��R;dBf�#
+{�b������j�[$Ե�I���ZFb]t�D�@-����O�#�[�vUSRQ�.9�y����y)&�|:(��� >�Wݯ�Yhb�"��s~����Yn7�$�,������s�7�@*����0���|�� Y��p��!�5L�Ң�wGg���p(�/��U�w�|CI��ѱ�0�˪4D��Gk��B�|j���,}	"� ��hz��Z�%�w.�0=I|����Z��	��bG��]������*a�B���I"�ؓ����v"2'��Y��7\�6���=�~*+�LY9,���X	5`�k����`P�U�������CΜOGٓ�~V���h�>�j�)��q�\�qv�Ю�{�v��1@++j_��CX1�3Sd	#B���@I����/������������Պ�Z��k��,}�uo`�:{�W�|
�Y��8:/��O:[8O��W7�ҦX(w�~�a��t,�m��%�l��Q'ۅ���/e����1mZ�C1;h�6���i`,�EQo�@��x��G6
��7)Bxq=6��`V|�d��T'`�K�o�*��;G��}��"�xrz1��	
�m4��.
=|o� ���!���⎗#Bt�XeM���}W��X�a����:g�]<�^�0��bKN��{#�_x�Ws9��,l� �U{O)q4�d����$W�	����ϫ�j4?>��n/��a��L��t���T�r�2f��Mb!�R�tU7�Վ*��e��@����	���QB�e�$T+� p Bz�: �ѭ�}�A�I��G��
f��C+eU�,�}4a�{��M!��>�ƾ��I~?+�����%U[���@�������R��v�b�4�ٯ򘯓�M��㍘;3|W���W������u���Z�d����w5���O��k�q,*��,�V3�JXn(����z1'��[��ˮ���Tw��#�	��1� Y`�%u,�������UCC�6Ag��!�`�g���s.-x!tHb������!��\I|b��kn�=8�ء�����\ؼv���2���x6�^neru�h�U6�H2?��p/��,U��Cx1{��ۛ�ڸ�d8/Dq���^�S-H|��x����j�����ݒ,���YO��@
�T?�t5t]`����\c��dQ�q�V\������2O����p�@qP���LS1bӨ�	5Y�!zA�^v�"𴏮�P��>b+
�����[�p\A}�ݙtʍi��a�h�fJ��4���K��n���ڬ�Raqt�������pu�Xx�qA���>��6�3���%Us��!�����;��X.���lA���3/�Y�Ѿ�/#�ӿ|k��h�+?�|���ھ��uGG��"u����|�Ya�?����q��nH��
"3H�EF�
;m�Ok�7�U���"4��������I���0����b�#�n_�Z���B���оVY[hk�$��h���,3�����߳��DMĹ�#��J���8���5r�5 ��)���J$u�d�l?�*�ʣ~�MW���>�|+�LUsV������3��p^��MFu�t��(��Q�$Z&:��[?�WL?�ӎ`�o��1��Wk�KZ'��ٻ�#	Ӵu��=��{+$Ƅ��Hd^wc֢3��
B�*��6�욉��\~	[m��j��X�p�⾿s�U���,������og
�LI�<*�u�e����7�ߥP�^#+����z�j��w�3�t$�I����mWPKX?A�&���ё+ZO
r��y�*�99^�-��fq�������1�!>�OA0Ib�U��iO>���mt6D�i�r_�!�QƤ���-\3ʏ�DJ~/oU~.���!��)��]��� tćwX=f�B�����I3*aI���i��
�p��lu_O��(�Ԣ�����kO�l�����;PPY���/܇�gM����Qɽ$H�UA�G�}<$=��G����\���=�뎰���5f�e�|b-I�7p]3���u_m6;�{,�h�(F�=�E����ߘ;^i��u訹�o�름��m�J9��%)�������m쿎3�S�?���ٖ4�����m,�X*�m^Z=~���q���Vځ��s�����҆-(=���x&l��r��k"�N�GNB�h�z'}���t�3wo�Y]����}D�	���`��6��m��ir��I���.M�%��zP�U�����Ƶ���d|���Y*����ux�:Y ��Z��Θ�f�;�M��4�y�P�u4K��g��Q�Qr�9sԖ���:�E����@j O��8��%dژ,�L}��a.��X��8v����,זic�o	�C�_�WmThYt�%���d[�s��;*���t����ۨAVh,��G �«��7lF!���z$~(�u0�+5�ǚN�b0�r��X,�K��v6�GK�Kt���X�Sd�Ny��Ά�[���h�2�:k���RB����^�hxF�6�H/��� �q]8C�Sl��g�xw0���ɰp�OA�b7@?������ǜ��׾��rI��o2� ��mb�
����^.�E�V�(�=h���ӄ�9:��C�����p��?�r����Q�-��{�0�m}6��y
��E���<�`�0ح�!��*�1gј�ǒ��)�V�S�x�����p3N�!��ہ�"�j����.�8�bi�ʢ����l,��ɗ�p��aw��C����R`�$X��#��A~`nW���PX��m�0�������:T�cTp���2�w�1��L�?X^�����q_g��@pv�Ū��$p�49��z�R\�[C��7翑��@Utzr�@%۫��� ��G�b��DtK�Ԏ/�=�t0�zP�^v϶�ר70�V��
/��%��no=*�N�g��F����aG��3K�^�����ȹp�` ���`$V}�)�v{��~.4;J����m���:d�>� �WV�'s[h\A���eV�4Im�}Cf�	��9\����N�z.:p�btu��(�{�q��CY��ӑ����/�T��in�؅������q��)�AZ�mE�15+��>�pS`�f-�𭂭�����C� �}��X?l§m��X�S2,�?ֻ���f��U!��O�<��{v�� ��?BV�Y��3Q�$����Ty� �z��(��/�$����CcR>D�����Y[��%�ו�&f��0��6U^��.�.���!(%\�]��8Q[`qn�d�}.\[��vL*�*��~p�*����Q�ب��]煾�Qq��T�_tm��Լ�=�ٰƭy�י˝,r�$z��=����%Ы�5��"b&~�e �
 �	(��C���S����إ������.�;�2aX��Q7�b�II� x/pR3.�[�3y��W��0��i4����Q�;�� fy����q��p����J�6C��j��n娝�^�~ֶh�g�/:�"�q�n�����Ğ���d|�K��k�"��&1o&T�����H�{�heظ��?N6F|�"����9imP�$Id��=�5U��t�@�~ZC��!*�m�E�Q��g��9Q)��J�dOiN8Y=:�#q�Vc_��E$�S����m��T{��x�4��ӿ)����R�4��2�9G��/LsT�d8];;��=�b��ڞ�*����&��G�fɎ���%�m�E�8k���9S�w���A���4(s�bt��gD�Kh��v�(���ݐ΃�߲�ξĜ<x�&�@�$۟�Ҙ��R��ӄ�Nձ�Z�Uܲ���_
��gr\>D�ˈ�"^[�F?�E����X�.��U�e ��������� J �f�;?l����y�-	��旗R�� ��Evy�2�$��F1���V2�5��c
<�c�zT���>dNU>�<�����Qk����H.��J#�~���?�
{�jV�\��V��̕�/�4;T0X���'o��_�H�W�|o�j�����l�vv��4����Ãү�����%�n6:�-G;�s^7}?���}�a����u^q���'Y���#
DQ����ؼ�]DEtN�N�����9Yw�}�T�z$ � {{��[�����j,`�\�5a�*��.t���>�w�L�&(���*�o䌯_����e�zl��øW����@�O��{�m����CC�*Iv���,�������Tq&N�rD��Гb��죻"��n[�����w�0P�5����^��( �o��ģ
!J��Jr͌Sy�,n���.���)��oIcO"��� l׍RER`?T2����FZ��]�B�,����"5��}�*N0���#�SDr��zH�k�q�+ �2D�1���L�+cd�>�VD�\{ڳ��O9�h��^�������J��8{�-k��R	�-�s���k�{[)&�t���B��ag��0?ƔkW�DS��o��1�V�(�M҄2�����be2P�5�h���?j)�%MO��[ӆ9�����ŵ+�H˃�f>�7B�Q$^�Au(�	؄W�VCu`����/q�z4�I1�+v=��E���W�j��˝��H�c���)Ր��`��҆N?;��|W�]�h���������-�T[]� ���N��j�:�2 '���PAx����j�kr�vI���Y�qg�	����V�糫�\�]��Û}��6.��1c|��y�b}�
G�ٕ#e�
,Qn�/X���ؔ�mW"�����^�O����I���w�����&����e;܈��x�����﯍�S]) vN�E���;�sۤ�<��L��=�#��żfcj�{�'`�Q&Ʃ�f������l!�'iƧtZ�ٷ��#������E�j%œ;�ͅ��
4}/�rO�#��<w�.Ƭ���{�T졙F�����ea�u�!���Hy%7�,#�,=��*fc����@�5b �����"!.R��IE[�(�(��)q<\;a�¶ i'5��y��x��)J �C{FΑz(H�_��G�Wۮ����Jq���^8�v�B>��	��\�>UβC�MIE�[�$uN�jϾL��n � �[񝰿O})y�V`h����d�����,��>,�X������~��7@&��,��.��1�V�kS��	���?t��:�xx�Ӵ`���X�����?����?V���Ax��x��u�+J�J(����[�H�y#���,(�~L�����L�CU+"�/y��;N�U��"7����2\���mh�_�����R�  	F�ȷ�y�؍��s9�4���"�2��6;"9�o�+v՚Ya�,2+�-�շ�G7�@�l8q��#y��,���ʿE�]���:�I�-~W���0���$c����6��2�{�z_��\ǿV�=�2g����W%1"�~�]�c�����lU�2������������T��}�RFp���hŝ8Kn�
�D�'�A�2s�#�J���%��~�́��6�J���\ �d��<X����_x��Nd�k�� ��B���]Ǒ�i˞��O�̥��9�ՇH�ܹ�`Oܗ�ړ��~�y%./L~چwǺA�k5D5��}����r:z�v<W\31�<�G�H
��d��0������P��
�����<8�Nk0#� ��G�<x!ojp
���]�n���ҭ#�Jd�?��K�𠱶nW����i�_zr���X� �ծΧf�}�Y��U�	*�L�#�0CCu�@����(����Iq�<4�ݝ��CZ��n{Q�,@���}���5���E�c6�zY���xR�mc�hd�B�$��U�{ٝ�䮗��Y����s-����1P'�x�ׂ���ժ;�&�d�w���Ԟy����R-;s�J��"��0�#-�C����3�_��֙�'Y�0�v�NIAE_DCfƸ\Z���ADU���g
I�<�o�P���uCUV��!<����y<X:0aK�^�x'���ve��-r���ľ%f,��x�g��������s�y��B_=��ьbd�}ݲt�$}�ۇRu��������e=��?��mOV��+���t��2��󊂯���0�9^�i�+�>�0�K��gI��K���ұX�2i�]�$vs��i��6	)��QlLI���P�?P#���sp�~v]���n��J�T?9���^�E��2G�ER���h:�8�?�	Ƹ�������u��U���>��垌�*�9�N�}v�-�%j��b�Mˤ�}��� �;�C�g	�"��w�	K踻��u?^wfo?r���ϝ������ ��B�e��^�8�6��0mED��z������ߔl^��=}�cF�M�FG� � =�i}���v�����^�}�����X"����ų.]˼�?dzU��<d۪��g�U�E�Y��ɓ-
`����m3����&�pFr��筂���N�t���|�n�b��֘�?1�3 `N
o�Q�����W�mk`���@U�����45��F%�e/�iAp�� �Q��_��4�[ÙȲ?3�F�!E�p����l�)E&����Ϧtk߇�8Z!*�f�냱��T�tgt$	���cfR��e<������vٹIL=�	i��!x^�1����k�ԣ�0��զ�E�v�aZO�l&�y��缱c��P�i5�/M[�������X���P�.���&��2���v�"�P)��<�i�t���z��jMf>�����K��*���]�E]�Q�Ts��