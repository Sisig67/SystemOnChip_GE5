��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj�o�v{'��p��z�ɉt��(=B���J���b�,���X!�c:��K��|屉�?�2SJB�oղ�?j��/'�]�
����k���~��}}e��X�!9���)���fO�Ǳ��ӭ�uZ�񂅘0���G�	��M��X�N<�������d�.�9#N.Ɛ�*F8����0���x�B�v��D>Z� ����{�N�V쑲Js�ϧ�{�(|��{���Nְ.�j
���-@�����v���5��僔�&6g��n��.xU�������`HH��Yu�Q= JB�`Xt���Z���4U���8�r���Fuc�cc����g�?wYi���P&�v��^����w]�����ӷ	1� �V��?���W��wc

0�:z��f؊7!��2%�2�Z�/�O�;�m�>v�"�&���;5&���"�1U�"~D��'���|@Qp�j�R�0sVW��d���a�hUf@�~	D>�(�Or�����(���L����SSw��r��r-�Nā@2c((�O�����*h�x��h���r�39B뾇|��}��)���&���:�0o��F��W�1Œ1������:��/�Q�~�O��vs2�YҌ[��I���-!0s��yq�'�3�U��t;�JOi�L�u4/���~W{'�P��B#
��sN�H_'h�ܙH?k�����d���[R�b��-�$&Cv���-~�[�d�,�ֱZ�F�h&]����]S�iq��Ҳd UH)˰cWK��$>����{��]69�W�����j��osp����S�b�.�q�B�f����� v)�X9��][Q���������66&;���6N�g����b���Ti\|{�:06�Yq=�%�"��а`�� �B��M�ϊ��8Q�;��z��
��K���V�K�����`U����\���m$`l;	FW���~hհ�w��FxGZ��,/\
�b�a|Dr�e�]�V B�Vv�!`2|>k}'`+t]1ޜ�G`�� G�Fh���y�!�儧��!]�h�pA����i�
��	��nw��XЎ^�ҙ}I�U�����r[�hm���bi�Ϥt4�N9;F�D�:���ԣ�c��)��T��,�#K?ܫ�:]ͼ="��"�=�"'<%��(�K�������VY���ɜ�
fq�!GH7Uz�m^	ݾ����u��Q�S���[A$�?q�,�jAiQ�0�P~��~x��.ǜ�pj�d��D�]�����yػ�ș'#@3N!.���V�Y�_`�+ox�E���s��ŝ6�x�g���7��5v�G���~�?��yָZs&�4k�痬#�;|6dے �#B,�H[`(OB�0N�5�M��L���1����u2��]����t��J���"��X]J�e��á)���]��s_v|'B�h�fۮ�%�b��E2��\�9����mBt�b�����̧}�h�x/��=�x:�}���6��q�5y�Gͬ|3�M�}���J���?�P ��&�'tl:��𿁆c)�`���m��K�`���JO������G����Q�lg�Dd�p���*�N�/\(Ad|��C��T%4�GWs������$�|R�?��L���V��s�W939$�)IV����Tt!y%���8�%�V��w��� ���u��ۑ�GN|�b�6���h�F$A͸е��U^��fƌ���^d��'��fr��g�u���?�\��ʽJ�A�J2�>��_S���S��#掁����>0*ꐺBs`�a��ɾ��M�s�Łؤg_O� Hhs������;�L	�9�f�����Ey�?Xz�N������ݸ���g��k?u-���dQ������`]uo�%7���_�w��;����*�O�?MyFM�y4a�I��W�f�.�pf�.�ja��h��.��/ueov��
 |i���qA�ٞ�k�Vfj<�K%~��LI2'��D+N�ly�-lV0�L����DJF��Z��s�x�|��r(F^{�w�$@YaH	t�2��?h�[�(�����EXGo����OE�G�:z�R�N�C�j��{���2��D�,����Z��bM¿	��ӧZv����Y�,����Z���9p����د�D�:1�=L��6��#�d���i	�_�����u5��y�px(��t;)�c]h�ne���CEl𹀆�r��&�X�ш`�*�q��iS�%�������SRns)1��R��f��B'�w�l�"_�'0e���ꑦ�2~��+݁���,�!Kٯ1& X�	&�G:�����*R笽R)����ޭ1�N:�v)���zIZ'�`�;Өw���"y�~m�,x�p��"�5o��[�ơ�'s�~`)��٘r���~b2��?r����]�A6w���߹�]F�P��,�1R��$�M�r��X�lɽ
<����8����>	\���J9���/�>-0`�1,p�J a<.�yXI��;2҆B:G�鑗�x@��8��ے_ԕ[�b�ʗs�����qՌ��t<2�l���Ы�c5%���AhԋE���dA&݉��i��5l���[�I���20�U��:EI�|��T��j���}1KY����]v�M����TՐ0|�*H�<�pǱ���P���?u��G�����dϨ�!s)��d�;�W�NUe����5��yyN�R�ޗ�v��'��q��ly�̳���P��������U�g��4���+�#�?pHo��ob��Z2BxWqZc������#�(��
3cć��@�n���5�`D՚��uUE�8~�vBx5�h?_�2��w�e�}���t߶�,�ak��|�'�9���P�'4�ۺ��Q�4���p��0j6G�V�}�׍D��>�=��	��!�	�o�@��Վ�ʮ[%�.SݓR�������ȵvJl��a��E�Ł�D�F��j:,0��c�ct�8V�Y@[�/j�g~m
lWC�ԛ�O�XH#7�{�IctSS�;-W�2|�p:�P �����U~[�0Oũ�/i���J>ݯ0��'��.r)�#�����k�Z87�?�A]�$r<=�������i^,�HkD��\ (�9�΋U����I"-�\�2�#�*�1�� �-(�J������%j{6�*���D��bJ��Ǹ�T����@��!�V�V5q!f+�P�";y�����e���I��[L1�2�[fs�)^tM��Xd��j�prC��TI6�l���re�cj�6!t�2H��ؑF��ο�����6o ܄�m��G�*���o�4�78b3�u�zJV����oJo�Q�o��~-��.�)$��gCL�[
 �!@����Ȏ��L�;�#�=kl��W��
�ޤ�z�����-��4i�$^`��"�+A�Q;�b���{'��	W�m�|e)��ib牎��.�YP2��IMf�.ߡ��L��-X��[�a���	^�I~��h����q�݄�W>�C�_J�໯!�$~�*��+#�Z=/i]�������w�BÂ��#b�,6`P�����y�ϢۙJ� 9n�1���(\��Q��jБz"#5��A [