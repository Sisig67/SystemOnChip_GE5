��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����P�^�Mqap)%t�?�&�Z�K�*���~O��in�ÇZ2���RG����R����k:�H����`�E�m��C�H��Ё�]]ѱO�UFH�Ꚑ�L
��"�0dF	�b5 �A��Q��+�	-�eD�4W!o�� �@G:�� ����Ͽ���˱z9-�n#��V�G~i�u^�L�������;�q�A�~��4�X�-�]Yl?/�Pa�����4ǱT|���G4'O;&�;�o�u���i~t��n���4-BǇ�aM�ݍa�ڗ_�bF�5�����
�s�c�<���w����\�_UN�΀'�D���+�qS�e-����@�\�By@÷�:K���F��W��MV�p'^���w}�#��
�VﱫIT����tL'c�>�F���b`(6$T�j�{���x>!���4f�R�;�'~>P�V���^�-x�v�:F�4�>I���Qn�0-68�jfb,:$�9>�X�y��?��vLr}p$?�Vw Q`h1���M;�qD� 8��_Cá�;!H���ޑ3p>g��;+F���گ$����`�͈��9D�Շ\����RrԎ j�JXږ?zу[@��;	��X�"���F���b:D��4��"�.�*�8��F����"K��rG�Q{�-M�ǡd�O�1	�9�^��қ˛�:d��>��1<�MaP���� ��a�0�j�\ ]�?r�v��œ�S|��A��ݔ`r��ʅ�R8I������-��@�(%!u셺Ħ1�3� ݿ)����>a_@M�2&o�Τoᇌ�3o��c����;�Q�U���{$:*zt�=����J�����ȇ!�S3-'��y���vC���3�!h�Q��O­�5\$6�14�9�2pҜ��v:nN�� k&�E��D.&��t>�
8��hJLz��R�ȅ�:Ѐ������j�D6B�s����i��4���Ţ|�I��6�ZPWy���h���ܪ`衑6;�Ɍ�G����-�=$�(��[�~^h��L��-��=����p�[�Nq�-��~ۢ"�\{u�י'�Ej#�2��p��&��z<�C��eFp�'xz�%؂�p�V�e�5MI��0Œ�?��Fk>n��y�ȹ3]����$��j(oAV��%�c� %�<r�
u��dOk�vʹ��Qh�d�s�@�i?���AB��O#b�Z4 �Tpo��&��p
�&Sbf>���xSIȿJ����g�1�3��-�@���r�r㪫�хG��--�� �ħ��<w�=�� y,����l�����X�/�Ñ�| `^s5��q�ȱ.���U��{��������0���Z�k	���׃1�y+A�i����7,��M��6�|9%3��+�';��)�E�@]�M<k�Ġ:�l�SK�k?���b�w1�"�EܥՃL�P9�B|�
PߏKx-������i[�9�2U���ꉤ�8��&Yq���
��W��`���D:e�|`����ždjH�Yt�Z��A��jT� ��
Q�u���*��sT�|��6�D��Rhv"L�4�=_����6~p��T�Q�B��B� �l�G�������&�l[PŅ2��͚W�p�>��~#p�N/��E��
�t�	TѺB�|PN�֑m��,��4Z�b�E s`�!^�h���n�h�f��(��F����[�1)�ά�єc8K� ���}��50�+��@���>^�Y�Ċ�[c��z/�$�C��#(�y8|��B�Uȁ�%��<csT�a�?���eZj���pJέ���h�C�~�I��q�]9)V=���;d.�evk�%�[CA�C��3�<������Btֲ;�
8�������W�� ݂ %\K�׿�>�qH{��gQ? ���� T�����((l|]s����ٍ�����|˄߽�V����O�2�x�4�LՅ�$��_��a�@��X4��2['��'��!�7�FS?d�ԫ;�1h�~]Bvg��V%�囄��1�cMZ!��|/��滵P�I��rO6�Np2�^��3 ����y2=�
�.np��U��ȼ岇,�����״��E _��~��[��)��I��u[.
�y�2 �ȏ#F��T��cr���}?��JO���I�����G#�<�,�=	졧f�'�� ��-��$/بN��̴��3(�"7Y
ʧ�t�4;N����A�-h���z_�d�
��@m�}�`����p K(�
�g��m>�oN5:�v�Q�X�V��X�[$�Y*��=�2����=sʽD�n���O����3� �@C��x��"�N5}��m�H�%�B��۝���µY�9A�S9��A��w3_�ɌQR�ʊx�_���%��
V[�ǀ��j���0m����%�%��
�fB��߾�g��A���Zd�1.R�����Posm���ڜT�C�����gpY�M^T�c��>S,�/��-pe��?."�pk~���������7z��ǜسw��5�O]Q���N�0��u�"���k�A�_^���0t�\	�y��+��/��
KmQ�Dͳ�h��^ױr��ܢՋ�re]�,�k�����osi�{�j���d�3�<+.L9�����!��7��mɣ{�⛢匉�EŸ�YD�t��_\���F�\�S"��m	�v	�ۮ�F�'��+��^-�;{�����'I��g�s(�^�dLŒ�������$�	oI�Unsm�Q��%�P�쉴ߚ���-��z���@�ێ�{K�X�6J��q���l8���W��Y;�r3O�SSW/V�]�mAhm���y%�P[�c���A��h�0TQ%���X���,�|>:*ա>�(�D�Y�>p��"I�S�����{/�)qa�H_��>�#&���5|blP�
���
���⻽`2����^���4M�aTK:aձ��y�a.���qKU9�ߩ���!����\5nr��p9�}Q����0��Y���5�Y��1s��к�>F�;[�L��+�A���򄩸Z.)��~u<!=����砨2�jM��P�K�?@hg�U�tJ�;��T�*_�Ң�qʮ��;n�^ya��'��GMf��q�����L��+���%ZK���'7�F��'5�t��G<*�XPψd(h���l�b���u����q��l�;��:4�e�T�(�#�^�=���;����Βgn�(ء]����wuk�Ո S�6���gZ �Jfa�Z�D�M�#� W8N=E�ö�f����^=9�����V��V�٦j»g32��{�)�m�&.2%�ґW��0�M`{[�)�����H�VuH�_Z�a����Z�-2��2�'�{
�y�㥄,C�����R�!�j�����: n}���&C�:�b�]��*�,��z:� ��hA�(�T�v0{iڍ����������a�I9Rp�u��W-���2���wz5;�"��Zjc�栁*	,��`iۮ�2+ޡ�p��A5B�:Ƽ�2�'� r��P�&��?��m϶D��AA���߯* ���<�WE�p�E�8�$L�w ��:,I��᥏�
��s�mF��vi�'��hJ��D�{a~�j��I=I��?XY�3SM���׻D�dCuM����aI?�ݛuп�G�-���HP�~/1�6K*��A]�b��+.M�;C]���������-UQ>�A^�]�(�N~uu��^�8��vg�,5�v�S��E���?��a���<��V��*J5 ��1ӛ0j,�+)�dR�����ƁS�}��nZ��A`�� v�R����^�a*��Ä=4��I�%��]T�[ܝm� ��e��\$�f60?� �6�N+B�l6�f�0UC(��K<n0�b�	ҿ�]�S��V��=�!��H��ϫ�RM�jH��i��E��P(!Y)�[�:�U�]6Ï,�m	�_�����F�mP��8p�9V})~i�w�T�P��WVDg���h�Vӵח�"����
��y8���kx�r��6�4��x�L1H��
᷁�����G8�K�r�9��Rf���@W5����)[�9'V`g�c#�>���*�Z{���O��0��
st[*��K�����bͷi��b�酠��t)Z��>0'���V�K`D�<�[�V��3^�#�y>i�2<ٹ\����IǑ�5�Lτ�N�dE�.}�/@`c�yD5��V^5X!��3&�̖������e���L���b�@6Fo:�o$�#����A���D���=.�O:����ѕ��aM�<E�y}�@�L����pkR�ڳ���j�$���������#1���]&��\I������L<��Xd^�f�_ ~]m�#S&@��zݓ؟���?;�o{C7��3���iEK��m+��*����bK���Vn����A�S�@_�V�ݟ)#n��1�'�B�!4c�I��V���i���b� �(]�!WꇷF�P ���l�����r����&��-�@C6���sT�Z�E|���O-�}a�J��u����Cs������V`�����C�\Dx䣍��H�Y��a�|��kXS�I��X�m+�Zp�ַ��4y�m�����.eR�4�]��E�L+?fl�x��9tg =���J������ގ�>b:GǕ�N��)N׆��A�ç��4�P��i�\.�w��H���4��K�!��}�>0i�9�l�gPndrk$[��`e�HG�MN���&◱kC6��;fe�g���^y�@��sk>]bZ`hη��3\��]�|�&�Z������~�u�ޣt���7��)��1^�;�-��ʕ�Z����-`$�D ;@5VuFƤ���3�%O��Ѣ
9��^��>+;��V����}����0�c���T%��J�'�j51�g�A���%�+����@�%#0pL�zr\�R 9Mv&�VA�E_aQ%in�ŵ�����d��(�F��vX���r��Z���K�'㵺}��7fT)2�*o8��0�X$
�?�&q	��^�%���E!C�5�9�n�?��
5�x�aK
�K6�H.ٽd�.1���Q�{�݇�Li�_� ŧ��'㈯�'X��/�V����:�N�i\�Q�X��k��
���@.p��-�<�5��Q:|�m�fW�F�S�8țL��,��$��%u� ��: �x�V�t>h"�^}T= ghhh��׻WP;c���n�\N�r�v�H�]�L,���Jy{��a��&'Sb��dP̋k�0g�z�i�z8�\���,Jo$���5���v.#ּ,��*wN��@���X��l�R�&�����2��߈ƀp���9������#?��*�?����jtl�cX�rm�:ԍ�X^p�*��|׹f�����7����w�*�����z�R��KE��ô^Їc��+��=$M=�EA�,TGj�Y4p�;m�s��C��[(��<#: ��B*yz���QQ�����ip����O�2)Z��*H�ԾR��n������iIQ�;i�N|K9'�1�K>�1��8�,=����(l
��8�{`�X��o�:��\~@�b��L��ON-�-��v��� �*�nt21�L�lyO���"�V�3��b�Ԁ��ӎ�o ��+�.��H��yt~=�����hf�_3���`���D85�� ��7
2�!������z�Gf�
k7�������~>w��)s��;����X�3.)�|�����]e�B��	����:�B�#>�� �î,#뼛�>���Έ�MY�S]!<O��0z���""ډve���-��~G�M��\)F�t)=c'�쮉�n�z�H�ǯ N7�,�<q�u�p/'.~���	sOڬ�s|vڲ�}U'�W��8�͹5�R�鳾@ģ6ܧ�BII}�W�n-c��4���q�`7��	���B`z�\�?ܬ�dM��z�e�7g/ƈ-č�`��&��a�z��B�����$��>��՗~��$�>�%���?��K{��xl�ѪW;�M�NxEoA��(��b��}�E�G�#�K����v3q�xO�ޮ�����9( �j���W�'������q4��!� ��8�<������6w@	wŴ��uʝP����ś�J���u����Kp�ubh�K�'.&ġ%�ض۾+	�
]yQ:l	�rj��K�J����u;���N�Kx��@�js�o��U$�,Ң�:ݙ�5�P;eA(~9L�-N�K�1��$gݵ�o[9z݆["�+mY�2QQ�T��7a��m�k-�<��9���,�-X�ٹ��>V�6Y?�N,u�v��N7�0�h�;�H��m�i`�W�IV�����M$���`ʼ��0�߀6���᭼= ��5D�f)ř��}�3���ӯn#a�Ej=[z��X˺;��bץe��TCc�6d�a��6���SO��ہ1���9��������3�])`�ȕi=�ĹQ�Ⱥ66��)�wl7�w���
��BV�u����#e���L<�b���L��YA�+�VM�	A��㫵�k�N�f=T�>�sW���T3��5�Ж��̰�	��Q�-�p�q�tut��dVm�,A
�v��%�u��EoC�8���b5Vغ(<���n>��Z��q��K���P��\A�n�{)sN��)^i���qC��F�:1�"Q���+��>5���y��nW