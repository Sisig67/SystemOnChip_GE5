��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%����!�rr/I���b2}���Vp��|̖�8��!��ވ=7���d�W��VfL����U	���S�>��E�s���O��Է���E��IZqGH��"�*z����m���T���/О5/b�Q����Ј(V(h����1���ʯi ]g�f"9��d��%�Κ��(�Q��A�8&��׍�% �ۋ57��֭m�CR����tJX��ai��Y��V�0Z�L>�y�?\���2�;�I��3�#�6��!��	ƀC0˴7���~�tH��]fj�+�p��;(3t��?��h�~m⣿P��Z!��EÜ؄]�j�I��_���G�	\�y"o ����&�S"̪M) z��$n�"����rt�O����%@$_mg2���7�"s��v����fբ/�_�k��Q�����>^���p�TuE_7/i��O��2o@������K4F*B_�Y��3�j�I�4�Pe;x/0� �#O!ǋ�C���2g��pG�x�֌H�nJ#��%��773Fj�	�Z��A�@eǃ�m�NbO����~�Yk���S|������[(���>��	޺6h�b9w��+�7xu\R���bd�������!?�w�S��r���^���C�ͤ�˜�"�B��$���
y��ً7�N���!,��7���d����!D^��d��0 ��mjh}�����Rx�"oD9f�l�G쌍J�*̤2;��C�� E���4��$͖�b�N���S�;�4y�Њ*��rH5nr�]�)j\�J}�Zp�R�1����|&�z3`Y��{�rMPu��� �.7F!�0E���_� խ�>@޸K��mpeAԼF��)�Þ	@Z��2�f��
�X}�OR8$T2�4�
(#��k�8�*M�����&�&5[;����.�0s�퇿~�۾}��H�|�-'�_����/����u�|�r������U5S�$���-�b�L���YP�����F��3�(���=�'����K��H[~�P�^;��p�t��a~tSI�O}���^ LO��^_}.S4v`���`m�d���+���z�'�k@G��}*6ꇳMǘ��0�T(�����iT�ȟ���C�{����A�X��O6?]���zn�XM��C��y��M�j�d#����S��ӿn3�|Yu����)*^���-�e�Q mo��x�J����=���7\6�V2��x������#��`̒�����\�~����$��u?�^uK��v� ks����M;�eS�t��;�.�տuVL��~�V�W�$l%t/iZV���&���WK�WD�Zр�v��#|esx����2qZfy�(���2���ͥ�|�N"���fh*V�E��U��� ����7� �!*Fy��Ȩ�G�[ rփ$�H(�wS�	�z�".�IJ~��uE��z�~$���~v�(~�fQ�Rй���c���Z!м&)�y��F��(�$�v����%�z���@P��u�tO��ɉ,|�T`7�k��/@[򌀖�񄐮�����S�a��3kշ�~�