��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj��_��� �@ka5�.���32�9�A��;B���No �m��[�a���F�IUr*�{[o#t���;!Lr�ܭ��8�����S)��a�� q�56I�������H�UX~+Ͳ�s�|M�����J����i�ur`�U�c�pK� �/xǈ��/�{�ׁ��fv�̸�Ӧ�C�͏��d�G�v��)���}Q�=v�g�3,tّx�粲T,��3E�<K,0f����?��7�t^?���&��<%Z+�sI�3�Hl�T��[�-b�:F'ڐ޷�q�N�@�J��̙,����+�ؠ��n��f��@���	)c'p��܇�fm��r�(F�/���bA�Y�cr�aլB9�3��fN����Ų�_B��~c���>[º���[�q��>�^��3�W�*�{P1�i|�vbP?��ncG���0�̳h�3j�r�Ok�[
d2�" C~�K�)��lZ�|"+���5�폲[�����G�Lm`�"����h.�(�<i��0tU��!ħ��a(�a�z����%=Ʌ"̡ta�s$.Q!䚲h�l�k�@�6���G ��IŰX'w�jd�.o~�kbӮ�[LUE�O2 ���YmxZ#oAOz�\ߋrÊ��C6*v~�d�J3xVb��0�#\�A�8E �Y܊��PsB�����C�yaf���OI6m`)W����U��@X��'����}2@�p�4�SOq���\�����H4�#;�n���+L�q��|Kͯ9�Q�I?�,:�I�Z]T`��X]WN8W�T�+����4�K��
"��" �O�1�	��9�u�cI�"ng�i�zH�Q�ͳ���A
VWpBw>��M��"g�(EE(K��-�_BBs�|���}�P�xC�H��^#�G��}}PT��yI�׌Bh�;ܼ2�i�������RP?���S��hɦ���:l�^���,�n6�-8�P'%��K�^�\
�5S�xC�l�U� 7U�	����B��� �ᝏѿ>H�WvC5&�%��n�]��O���bFl:��q\�`��������Q�RFx�-��eܦ�I�v]�Y6�&w0}�6����)�i-K����Q*�I*�<����8����L���ÊKV�\8�\�D{��"�̿1��&������h[P;������.G�Xf����c~��EY�:������gɘ���%�q�V��bلN���1}��(��X���R��\�bܳ�-t7�!��C����Uql`�ߑ����Z����4����].ߤ�C��D�Q"�BO��\U>�̮�;��}
�'���$�Ӥʫ1�A~��jH����*^iT����|��G���(FjG��������4��u�B)�1�����D{�t��s@�h�řY����!ʮ�á�E,��_��c�=���9�U�����6�l�ݾM4�xN�<RH���DH��S�L��zmN�AX��7�G��r�Y��=pak �1)�y�CpPde�*����f�u��C
"�4A�i<����_D+ &�}�yS���ߡw��^��k*2�2�G�l�I�x{��Op��7G�z���j�D�t��fm�%�7Y�ye�1k�Β�&	 ѝB�{Ie��W��`�j-������m�xr�JU(_�	�7���G�,0��Z�=L!����/�����r�1��W��L���{��m�#_�"�]�97�fm:>��m"Ok\��_�{����h�w*Q�����,-���2+{Y\A��k�77�ȍu���5�	��t�^��v��i��x�)�q�{*�ǦR�q���Cq	�͌ _j�]p�yF�`<ϔ.: �X����^���Kev��6�!�!��g�R�3��җFM3@Q���A�8b�؛�4�}���N�Z�.;p�T
�������ɂ�{9V��jz9��h�.�����R�����u�Yƥuy��@�l͠����ԣ�T��/b!y3���,Gr)�[F�R�خ��8��93�����Z@������Rh��Bʖ����g��.I;�i�k�;����:�y���q(�EL����p� �:�3_�n�MX�<>����ٴ�t_a���܁� ;��='�e�WQ���ȁI�O�����q�eO���0���V")�x����וbv5���!�Jl�B��ĻQJ�>���}c�0���P�!��"�����+=O&<o�����<g7Mt�"�	u���C�����EV=�lyc��^-�#������7$�����������2�`W�7nH�=�].�F�^��������v;�W:5-��'Vm2����ŋ��_�w!�����O��m�M����py�:��4���Y����Jd�eݔqBjz.Z�t��R����2!`Ҷ���z�{�cl�!�u1���nA֘䷲��s�Ǩ]@v�K�_��:��H�G/� �{� +j�`{e-�d��4���p��Iz����'�����H�YƱk�fg��O�笙΋kV������ ��?vP�fF�-�h�b�hO�c�K�����%�;'�p7M���L�&.d����<�@EB��,z� =�rb	�k=;|��~�K ���q�͹��[�ʈ��6�M#�S=s+h���c	������c�C�?4`��.��4�7U�往mfCq�QR�e�\�]�Eri$n�MWw^����7�v }3�,�oCצ���py��b�n�bw�ћX���Aw�il�T*��8{�N��T��?ՍN:@��_F���j�!d:��)Mr��{���@��	��^o�/d��Y���>貂u�ū�׶0��mK�������MSo�D A�f��a낀�����t�WثL���V:�W���6������]6�H��M�2 �	����p۳��P��(���T�ggⵟARŉr<���)����Ń�v^%�8�ǫ<P
�ILr��E�[���^�w�y8:J���@���T��r�D�jwЗ�mߥ�D��$(K�>l*fng~�ܘp��,�p%�t�E�~q��">սC.�`�Pt��B	R2�J��r=1���}�%d⺑��I�r̆욧�N�H�:��/-$S ��g��z��}�^?B-$LЅ��3�<�ޡ���f�-�$a�n�LڅZ����[�Bc�}��U
-�CSV| Ή�#c1�F��^��4��il�O�Y������`@M����G��j�+/`�iX-�[~���74ML�5�x�����p�q j�\����U��`J�H�*�@e RUN�E���H���]D�;�&�3lg�/�{���щ��U����8>u�����M [M�P6���A�IMHc�I�� /�ao_i%]B?&\���9�y3�<��ۅ�(1}�n9
ĥ(���-Nx�����EE�v�����l'�����*م������ʯ�]>M��V*��N�I�V*���5>�۠we�����'���ۅl=��0�}�p��?���t+@1v���d��N��ֲ���W;��M3�X4���L�Z�O��;������T��d'�]_�5��d���qc/ߘzCT�S陝,��t�@@uu�2���c������pI҆�w~�L֬�<e�E�Q�[`�/�4c�:��'nP�ъ^��@k�����I[��c^^���؁Q����ߴg畠���囙ƹ%^��!�����{��JQ�*A7�eI��dn�G���z��Ln��9ڛ�-�%Vy��j�Z)��x�fe����U��r�����b��t��ޅ�0�RX�+Kn�� %[��)o�?�����ćA��<����t�9�������<�,�і��/z]oCIo��]��z��S'/�x	ok��&�~E��xhȩ���T���C6��>jW
�`�&�w�
5�B��$<�Ҵ����9�Q[y�� ��6�6I1��G���^`��tk0�JX&����Y��*㢪��D Й����3�w�N��%����j(����i[�KA]����&ǿ
�<�vW��_o)���Ci�Qr��	o�x+Sv��`b��t�x;�n��e��b�
�|��*�B�-�E=�qL��l�5L!��\#����`x��aZ��z�0kC'
�jmܰ��N,�0��ID識�V�g�U��4 �z��ٿ����V�Q�x��y&��vq�4§X.�$�'�`��&��5m��x4 U-�=�?��s���y+�»מ����^rՕ��Lf$��L@6���K��	�D9Ά�;p��V�Cq1^��4�&�P[�����K�¶lӡ�s	C���W�C���!%գt	8\L���S��8O�n����ݏǭe���"� �b1�=�_"�K&")��������M�^c��@D*x4a�]`b�����JA��:�������m<)袥�ſ���߄�)ʤ{l�3�٧� ��-rپ�i[\�j�'Θ��»O�������z�'�p���7V�Г�RK_x�B�А���P��~�W�u�.����,\���=�"Y�3�@Ė���0"��=2�6��*[\*�5�8ɾ�� /I�5bߴ+ �����(�,O�K��Y�~�x�{�R�f���uĶ섩X�A����~ퟪ�z/{���TcTdk����^�l>��E��F�+�gTK�c�q��e�o�:�C���u$%���SeI���."h͜>����ER)���Tn�T�a�����@�/.[p�rEFr��x��|ަ�V����%~�d����W�b*& (63�%V����3�Ɖ�cխ+�!��U�vO׿�����M���F'|��>;��J7�1�`U�c�G0�J�࿨snw�"�vQ���;��gA��r���z)ɢϑ�=�Ccb��T��MtV�߫_��^�* �"ĩ�ke�j�d`H.H0���z��t�@�~fphg+��!�J�f��I�@q��9s^���U5J���HM�X�;)�q�@�bvf	��2��˗��L���^���b)�~fOh��5&L��[��t �k��@R���~�a0?A�aL�T^�`�3�������z�@H�S�U�
�����2���,c���s���h&��M�m%�H����n� Gj����� =i#�toI�_-<��,�I�5EI�ѓ���[%����iuhSz�v�/B�|j䷎)4�E��|=� t���f:�q��ݖ�.�8?'(LE��1���H&���yRhe�Q��ς���{��+��B��bf*d䃲Y��H<Z��t G.5�q�p܊���b�y���+jT�4���_.{�" H/���Qm�Pܿ����]WcEa���)�2�C���������߱�d��AA�e	�13Ee��>�7-/�$�se=L>�f	G�nz�:-@`�
����.�T��v��g&�h֭�OP).��=Ϲ���'�=4'W5�}(��/���v�<)�'�֡���u4����&��f�ǲ�̫�~^�7�l#w8��n�IkJ(W�6�HZ��ܡ�b��%��:�s"ݦ��O��p�cj�0 *$����h�
%�Y��SR꺳]8��4|N�_���rٔ�w�#G�����e��Y� f��H�ґ��څ�s�E2��$��uUG�LS�?�@߯m�w?���!��b�n#sD�0��J=��hF��o>�f��Q��k�ilxʲl���h"%U�{���5|�q��,��]��*�G����&L���+�-����X��13��l��$ґ�h\+W:�!G [m ge�������.�>����{��X����4B�f��ر�Z x��xi�E� ����;xGጶn`�'�5��%{�bh�BV�X����a_9�T�E�e��z�|����t��g��W���eX}(���ʺ��)�c�/Z�A`�8,e��5:⚘�_���.ن:�r��H������ɴͯp��'~&h�ƀ����=X��Z��+BU	���e����-�ה�aC��"�7��I�ڹ�jï>�sgh���Z�4�o��VJq��qyeHJz+�uK	�$��	
۴�ƫ-�\ϸ�r�򶫙++7�U>F�9P�=���R�4WnPf�ׯK[!��4��(���y�s=��ۗ��%z��������ͅ�V�#:���?oQ�k�޴�����p����E&}ڂ��"��<#�rA0w��.�����-VǊM���t���0��;�W�,�"E��:��0&'�"�pC�p��A��8=t�l�s�1��c/��sĶ��[7��B�I��_��&84T���jL��Oɞǉ���LH?E�m��q�\/�D�IS�5��jE��}�-�$�
uՎ�.i�P�W*
�L�I)^p���޷i��R��M4y�A��'۽9� ��D��~4g���Y�/z�b*�4�R��Q�8\�v^ z��z
��O�����N�p\��j�e��kL�5Ɋc^�HN	,�E�� ��Y(�>EVL+���~�1^�:Th�}��?����T9u�ᮩ�/H��� �77/�J�{
��dh�ݼ�Kx�=Ŗ��L�����sk�]�=gx�&�����of�;�.$�W�f��7�;#�P8�୽�S�iA�m���~��zdE>`{�s;�}������7p����򄤰����[z`)��I8.��Ay��k�f?���hѐi4 ����(�l�~�S��N���5�U���M���<�B̠bu5��F�7�6�R�1����)�zͿ�A�S�}�f��5���8�?�@�V������<�T�I<�t�V��."9�'ժ��6l�r�/�m� �֏�dm{6�����3s[yȎ�	�s��5�њΛ�7�s ��/w�$"-���v�AO�YN�Ұ�̽��v<�C���\��j�W�a�1����Bp��Z��Vnm�����"w�!��K�'�> �i���o� �H�4(�`�ۀ�b�;߈'�f��Q:[����I��I#i��c���H���>��Qf������P�S�1���+66���O�b�L�ҿ���b��S�T/�>G�.�m�K##g~i������#(��]����bK�yO[$PXE4^�A���E��R!K�-�L�;��򭝻]��Lfy�\�
p;��`�&��:[�:�4:�1�ҎЧ����4j�����#�_0����`h��m�������\J_���ӝf.|ٰ�(h���oW:���px�ahʔ��c�����ާ��CJ�2�OY��t���<�DB��U�i=�����q���u�O�T;dZ��|�_p����S�.�%�56	�V��an�%�c$ځ��:�E\����9�vr�47S� `�²�3�Á��8� J<o��Ʃ�N�O�%	����VV
��9@e�4�\��VD��I��B�=}ڳm�#��L��h�1IT�	�T5~�X(���
�	�dl$#i��U�f|V3���a,)p��ZBw[��w�N�$�H/��Wjf�J��'͒;iʄb.�ؼ���v�o�k��%����n�UX��,�?�G�ă�	$�/R�˕�����;	_|��bj&�6���&�
�g��6����~��K��5�������p��e%�9j���4�vZX�%�昘���+r�`r����P�"`��H�x�늏�C�\_���N�mC�`s�:�����d��T<�XF�d(�C1���TڭZ�VGzrK2']. ��eL)=�������C�b�5M�ga�&��S؁X�n��{b�]�h���QƯ\T��F��S��6��̈́�L1(a�h��ެx��˒��O��3����{�-��@g�<�� �v�	R����T��!��NX���i��3��n��������}:�T|����%���AcW� ����,Ezt$ߨ�	o��ӎ���u��Bdn���ǌ�.�� � Į���p��3kHi�2d�[~C"X�H�,���Kw'�s�`<�A���wؔw �QWw���JO�Я9�P���rG�Pi��r/�o�4?̺�8�kG�I{jtዥ����)��O��m�C���EͰ~����ө��4���TlIG��h)�F��ej��\��#c�Pp6Z��N�,n߮�E�Aal0�R-f��Ƕ6܊u���0��5}b��Ќ}٘�S�Y��t�R�3Fc�H��#�T<Su4���JI������� e���YF��A�Y�!�ʦc����J�f�QD�f�ib��r��VGU������ԱcZF 	����f�.��XBlLl�������{�u�5�����z����5��hp�LZ�u�إ C����?R��r�!��)��&��.�g
�w7:p)Y0��wY���0��b����4o� C�r��Ԡ+Xf_������f�?�$����z,��y#<+�_���yT�u<��F�I���Ø��6sA���t�
�ٛ���e�����6m�\p�?�����Y���{����M.��LWD��ͺ�;:%i���
[AN�Iljk�Д �J��l9���%��{�)m�ɴ���_�̐N,j���]�_6��� ��\�aL�D����X�3ۂZ*���r�t���kx�C<���{��N��"����\�y����A-%?�&�ۢK�6K�������\���=�ц���t���}���C��c(�D�t1k�����jC�~&c�H�N�4�^U�����I������\{�����"���<`_^G�MI��'����	�>�y�;;=S�r��kl�<<�g����3�M�[r��b	��N@�6\S>���ĕ�'�o��>tR&d�Y��Dԅ�8!G�`����-���E����{c"��<�aR�5�����|��]�TM׷ N:������}��� d�}ROb�e9��#��	��G�0e��NY6�N`ǎo�[��K���	��U=�DJ�z���}?g�g)r��/�j���&K�c�&k�5&�t!�G���Փ������y)����~���q�� ���e��L��F�]	��<M�:R���D�Ȍ<����v��*+�K|�HV�6�TQ*����V�u���~�����ݻR�#2��)��&���L�l*����[k�v9|��f�Pe�����W���]źMt�����Q,.����\1b�<�����Z�"�A#bD�1���4R��뛂���B��D��*����5�;WD�RF�~��X�=ε�<���a}Ck2����G������)���Qi6�ŮSa�
jBT�s��m���g�������_�m.��ݢ�(��?�ܣV|�r������U�~��JK����<đJEI��ȴ��U�!���_4����W��:� ��zmL�A���8��l5\NxU��2>1�a���Qh�!2h��6:��BM��{ ��hB��`��5f�^��0?TǑ�}��>)YG�߂�G����@�E�	��;����_� >�"�GB����b�*�GN�Ua�+M?�n�,���B����M�Y����QA��a�d�`��d��s6��[O��)@ DT��6���!p��XQw�@g5��+�ehvVøf�d}�#�Zb�H�R}E�;{&�i�6pd���G�F�Niy���,��ϩ��M��f�&�O��9M��ۏ���@��+%{�(��H���3];F�'Q��v������4m�~7���f���NH�ږ��V��>�C�o���bXyx%c
3��(g$M�cqU��X�ݠļ�㴚7�v�/�O����[V �\�-�^�:�v�+Pu����j�b+J�F2�K����pPz�q�x���7ףg�(�8��0��{0��YT�B-���	D��􇺟u6�t��&M�Ʉʄ�]=����Η� BE,���QFZ�:A��J��/�M6�V�ѝ�j�,m�`��7�c�FO���v �����5�p>֔ Ҷ�{	�؍}xէn4C�*�Mmc�`�$˗��͕p��"������%SNS���L��W��u�����?�Ҷ�����7�<��!��p�?ǾE���e3��.�+ݝ
/��ӆݕ��&��|Д^ڄL�FWi�Owx��[e(EI���_O�r@L�չ$.$gʙӉ[��C2郸�bf�`@dN�E8$��6��eջ�y��:R2ʴ��I��ݠ�}~b�
�΋�@�kt�������J���ޥ	���রz�64��^��
��y�F�r[.)�?Y�RK2R;�h�������iH[� �g$O>z�}�U���"�f�ʁ�.L0^:Su���rw�;NЖY�b�<��A��RBP�;n�G�p+��P��L#�~�xc�=��S6=7bJ���4']���y=z`�L��K�(T:6�����ߚ`�@0��/T>5�J�iF.ޅY�k���,���q!������ Tj��B���$Vb�-rC*^mHo�*����*�;{�������-vy;�ƾ�e<]�"d�5����q�'q�AcM�$;���,w��^��6��u��0xo���|�7Ƶj�Q���I�c��e�А~>BWnkY��B+B����eR&�s�c+�\�d�Uu�`#aQ�f
�!��y�)%���n����@z�2��IA?h-�+�e���m��N� ��6*~���;���/�@ȑ���f����G<ǮuQ��_���^U}���%��c�%��P����̹1�5��{*ּ���Oyx��&?t��=-<V�
�U���u):ZY�-dXt����ww��Z�e$����q���.Y���Er���G&t��juף�8t��E���O�	k�e�x2V�vtf5�\=�X�r_���eA�Qe�}�h�8�_č�������صHW�e�8c7�zX+�Q_���m�<�����H�ϱq~�R��<�f�.~K(y8���z�*�i�J@��ꈥ��o['xQ�"�;	�.x����Lz��h^E'��Z��*�k[�j?[<&V� ���o%������ (`�q�䟍��NnV]|�w}!s�kY7M;6jd�wh<� �F[�����%����	Ŷn??? �ߦC��up�[aw���W��G�M\/�*�	����)��5[:���[�"ab�&�VPi�/P�<���x�O�{A��"�x�U2�.�}ڹ�9i���|L�'{9ػ�Bi��1$:�����e�[����3A��w2ih���y[:5������L�zw�f��F�9�oZ3j�~��V�]�٨,��$�US=���֌��a���%�e����j������Q>�9�ٔ��
��2�2�;s����7j���0o4��-D��G<�Q:q� �h B��ʺ���	�]�X��?�a@��@��c�SɁ��Y�C��1��go �0(<��Bq|����p.os(2��CܒQ��/K�o���#�p��N����
 K��=����1%�y^�ȭ��n��m�O��B��p3��X(S�Z2Q��ASpäE��J����g�p�]��s�=bc�|��������c:\_q�ts���-R���1�_X5TY-'�f[V;�6.�'���2���'�T��?!�Wh�E���������1��kV�g�(���	�K�?K6����<2��=D��V>����`é!tU��g����i�(�v^d3�d��9�������Fҳ&�* qWgık��[��N���(�HI4y�,�|"Pz4g�]LU��Z��Z�,gjq-*�Xe�
��o.���s�N��=Yē�v��|�<�����K!��LUJ:nqL�"Ƀ3��؈��
����Y��2�j�8+q��#I:�;)�՘?_Xh�e�Q,��NX>��Wn�[u�cW�j�D*rc��0S9��h�I���.���viJZ�P.�h~�W@i�$AW?�GjL4�/Q-[���&]Z�����dige���-���dY���ls��䃖-	)����|ʻ�P���e���/3�"�n~��T�j'��PC�	xڑ�����S僃��˲`Ԫ�l6�]���ȋ�_�ƿ�O�,~ҩ�I�0��n��$��+��6ɲ��E�^F6v ��҇����'L�PCw)�V9������AU):��R�.����˚n2o�[�Lԙ�ee��{�s�)��60}mx�μ���j�X젯I�L�)	����X�;��՚���q�V� �6@MM�BCP6� ���!����>�9}�	���>(�ۓK۬�'�6N��}y�����b�G��Ž�����E�j�")a2]rK0}Ð3�����<t�R	i@#���e�n�iK|���sCq�1�]��]���iO�ƃW^�
h}��,X����qwy�5��Bg6
�E��nc#������lWF��o��p�� ����N�xSdB���t�� �YG��m���D�rml�߄$I��Ig��:���,&Jv��+*���4ߘNQU���[`��E�|�"Wֿ��e���3�$e2�Ω�z
s�t �������S���$��(������[�:p�ڛ��e*��N�ɇ�V`mq�(K��n�o���wȼ��L9Jf�`t�T��y�Y����%0v�����`D��3����4��{����0bءL��ț�+:��G:�'F��q+�U0X��?Q5���FN��8�r� 3�]���g{�k;�2�.Y0�C��t)i�~�)������fU��j�O��q10EP�~���.`ɐ��s�����w�R��J�[�)���RV�eә��J��]'~ǋ���,�Z��q_'y�Ɏ��}I�Ty���|�UR���q`��@׉���m_{P�0��gI���VX�ikRޯ�F��.�"6���ID]�gVg�<b� ۅg����w���Bʖ[oXs�0ӳ_v�l���|�#���B{8��C�0_\H��{�{C�3�LF� �GS�Y[�"�qˉ�z�=�g�+��(x+�!U��j�O�1��뀥���#�VW*���oj0q5On��I���|k5�=~�S��Ɖ�॓\�ٳt�)���M�aw�6.3(���r�hSU����#�;�IT���N`�ª����	��qY���o����r�����b�� T|�V㑕{�I���by-���B�b����M���/?U�PK�1&��
5n_�~ׂ�1
��]|�c��<�e��b _i[��-��T�d���(Z����8�@�F8�_�jg-,��v�C��f����^����S�sdJd($�gt�M�=��vd�=�+B��$�Rtؖ�H|w*@#�V@�����^����`�)�
-�&�R(����ˤM^�3.��Gٯ���yip���dLA�?���[�3�}��u��Jp���~�Ɣj�� �$I��������� �"Z���n�2:4�2�xc>����P$�\������� �0��W8�n���a�!��n8��Џ;B��C�!�ȐV$�d�QI�Z���#�L ղr�6Fg8�n��I�mu	�H�Cb7jkǭ�Np�0/H����.g[��C�W-:ܥ�:ȁ�����w�$���UX�_EHm�.���v�r�ʫ�'���!��!x�J-�+�����)�)������<��f羦s�r�Dc��_��u]a��$��!�C���d�"+D&<J�DL���~8w1�(-Y��7�d�QE1�"#���9o=
_J��Tн��ty[i���7���sh3؄&��/��Mpc�	�bcF�O$ �u�d(-�9�U�C+�ʾk�i"R�zIRH��QL�*�����8����K�)��EuS�g�\ǡu���p�~��J+�`�� C��d�Ep��?"9}��d��uǒ4�`�)� ���
��`�V�PY-Ҩϕ")����DU?#B�o B��X��,�y�QeZ{�4�d	��t]|�#O	JƜpѤb(j�B�+[opIE
��2�Jie5/,=�8p��+\�8�$<3�d;[t;��L.9���sr��a��O�)@ؗ3�R�|j��R?�q=�P�-_���u/�u0LtL�(Ô��S-�G�Yj���政^Ҿ3��� ,�R�����Ji��W���%q�(b����D֙�OS��*�K�Z��Iљ�,�
�����c{I�ҜE[�ϩh ��v���7~Ŕ��,	���	�$�1H�8e��q��T�d���i���\�'|�f#�
�Bg��幛1���,��r���U{x�r,A���љM>��L��YB��e�fK\E�h9U����$85����6�K����z�<����`r
?͎�,�,�*�w��a@\`8L9��uC���ͼ|+6�	��Ln'�B�z^�3�f��x���"wN��P�×�x�:�`�5�2Z����.����v,��|X�J�����X�T�"��ey���{@�Z�(ޥ�'��	��[�a�q�fb`��ұC����DF���#N	��ı���`or�H�XÀ���:O�
��{Va���Q	vwg�~���޿?�zA�@y�׺*���!̂8��6�jR�xCB���P�1.�ĉ��	� ��g�b��5-�O��Y�wUI�n*�8d�'5��+a��U5-e���2RW����<�������	�K�w M͍����:���Kr�z���P~M�*�­<�I���$4��(�򐷐ԼhU������9H�_*%T��^<E4��)qs^��ZkW�Ε�>�'�D���	|{��"�~������D��ľ���O��ΦPh�'j=Ož�#�T̡y"x��H*�0�-�ބ�FH��*j?���� �|AxYV탩v(У4��}�PP$C �a��b�t݁�K�9g1H^8q�TNs��b��.����m��Cp �4���=�x5����=K�������P�7|B��P�Y�� ��rǣ�O�t����q����ى�,��1���;pwR���"��Kޑ�zR!慲^���M�Q�R�?KQd�3nN�̮��Ādi��i��o��z��ےG����p/� ag:����8FF`��t2殳����V��� �Q�be�CK�">Ox	x1�
�"Tnd1��GF 8y�o��辺왰���P�ϊ��5]~/3����_��!PG��Y����-κ��[�$�����*��AMj���--�Y��U��4=��(�}�O���2G̖��ra�l�W�!Q��{Pn���$��>�aW'�j��=O����Hn!��A��jW3.�N����+�b��������=��~H�S�04���>���K#w�,F�	+ b�$���V�1�^3X��N7rO�^�Իw-il�	�^�x7
gw� �����q"�v_ЈtJ�h/yɹ�S~�Z%�I�����=풟��G���6p��ye����(�x&�)?�Q1�n��ȗ�Ms��A��+�i��b{�|b�4��y<~�.�m���@�<�	����r�z|�-���"�kE1xgk����ѓ�_T�����פ���a�p�/j�t4e��Ip?������=$N-��;~N�ʶS�U���EX� �B��-�!H�,2�zaZ��RyU��o#x
�}�����*�≢�=�7$����<%��oV��!�[2��>>�
B��.�I��ɧx��L���J��X�F�?��B��_
A�Ҭk������������?(6�����D��J����u�m���us�K!�����H�����j�R�2t%u{�V��4��h��2�[ȶRȅ�`�?= R�;����.C�o�s+�\��&����v��܉������4�~!�x��V�vHe��y��W4lԕ+� �Њ���A��](]'Jyr!��ǵ����*�ۜ��y��ʳ�Zw�9�Џ8���!�����+�v��d+t��2���O~6�5�U�`�,��x/4K=�G�Ơ��Y�D�!V�u7�g�i���Gc�\O�P�=�?n�����o[�a\5OU?j��Rj-B��9[�M�?f#��r��9�v]�גD~���[�!�.�I���F��
�^�/P����~��{�����J�/_ �R����==���"�w�a�N��i)�����\Z<+r�}͑u�d&#�3���6
��3)S��C��M��+ع�=xh`:�l�Qt4PU�Z�0H���Icx�l��C�M �7@Z_�3i�K�8�����RԚ���Z䗔�u�fZZ���hlf�*N�U>J"�,Sl<��S��-%�7���8k�hU!N�@�C�4�e��w�My��{%`\ʔrcK[�L_u�#�i�kȌ����Yz��?r�>�f�X �\9( 9O� �ċ��܏�1���M1_&f(W�E�L�m���%n�go����XW��� �D���R;D�:�	�#8O��
�GN�''�[�)�d`g��#�H06�Gt E%�J�!�x\o���{���ݥ���d2y�g�]
��:��uD5O�i�OH��'ۙ��� 긍��6�kY2�|�$�{_�Ф��ݢ/����#m����!�%��FD�� e���m�ԥTe]R��G=�卅vؐj�و������Ǣ��<ք� _}��=?j���y�h�b�,�融�����.'�n��94�����o@b�G����bR���`�3���_�Srd�P�@x��=��������`�3z�{�6<X\],2Gh��eC��Y�cG�b{��#���#�fFj��f���D�ձ�!+~T����u�w1k�|\��0��X���f�-����:��Cer��(6�7Nt��0/ۺn)1� �kZ�|��Z;(O�A�
�H�v���ݬO*Z9���0��Z=�i�p;��8&4��I\h�BeY���cT��
����Ql�zЖ���w�Z�T�8�Y:trp>�i�ѫf@�mJ�rx߿8r0FCQg������WM���D�ZO���> v=2(yN�w�u�������d�?P�A�V�urk���qe>�
�e?�Ws�ť(-���É=�ʺ��>Nڙ7f��;��{���e��g0~+/h�}�E�2w-���Ht!ۢ�6Ol �u:����Mq����P,��3q��}ߐ�w��8�ϯ�$�[�Y ��;%�����wx��q����]���m�2�/�/X����|e�,�GTq�`��C_��͎w�찌�Pq�"m����$"<�Г���(�%Y}f$���2|��o��)��Hd;X?�nY9k��϶A��ʹɯ�7��ܮ#`f�e[�|c�N��Z�I�}L�t��dGHp������'D��T͑6/yo�s��9a�ޖ�|B���>�bO�	TE��⡐�ZK*�8��T��VF��/�*�%��$`k�����!ǈ|Y�ڂ}��!x���\mH��ӱ��,��G_>Ւ���}�a��#�4�Kb���/0����ZmȢ��O�.�Q����e�Y�g���H�Ƚ���Z)���/�C���2��飃�lp=G�&�oSȲo%�MPR��uު�%�Uj���m��}�Μ��e�H���V�d�	��>0����:���T�Ŧ�(	��7���۞�^��w�{#S�h_*��w q��O��X���>G�$=��������
�D��KK�0i��ѿ8�<���
�xڨ������k�S�]�C��(��I�"��"���5e���֮\���!v���]��� �mKCI��-�l�C�$/��^��ߟ덅�'�ũ^hu��=���;�%�¤���0L����wVo�U�r�A\W��\�|�D����gw������hq�
�7���Hbd�N����(]5��˗�ߌA��Ԯ�
�� �A.������`ia��	9~��D�3�íFrp���A�!��s�!��7-0E�u�2��2��-���꠶��0��'����5�E�"��Z#��*����܈���铴���[��9�SI˩e�Ƹ�d���0��t%q5{��۟���Pi#�Ư����[y�2*�����1��-�mdUvc����-�E�ϻ���J�uM�� <M?�����å�3�M�=�rb�
�o��Gr*R,�{Z���"�Q�%�fʔ�u���c���^��p<m]45ƻ���LԵs� F'���-uX>M�ҥ���:��Na� ���[�+'jv�[��$����`��:�~�?���XQx�
f�dKe��QS�T�f����Œ�a-'cu�"<A�:��t�t��9�yŇM��W��&!���F��
�N�W!�?�ma��FuT�c]��A,�|U+�Y�W��+�3P�yONNu���Ơ�V�<o<�I�Vګ�]?��*U 3KP�_�?֩(������nt��6�J<���ua�O+�܉������M2%�6�Z%.��o���ܐ0nL��Ы�
�|�#�C�.̹�z��9��$�k-����� v�8������#������9cV�9�+ZЈu��rEw�Y?U���-FP�=*�ٲCA��u; ��]��dbٻ��l���>
����
�
�YDy���������ː䆩��=`ɚ�P6{S����]��Xf����ó�5=�5���������Y�*�g�d1�*c)�+��]�$�.���?�ls��o�ӅH�[���/J�����TM�f���6�F����r��mPw�]30����҂x$��S@��+��42
�OM ��ϡn�=�/�Z��O��}(CR��b]6�8Ռ�n0C=�\u�b��?�w�O����q�}S�D���}�Mb�� !�=6wXH�ӣݜ�cC�;NYO��@Y^IXSV7I����Q;쎟;��V'x����`�罸RTqs���!�8�|��6n):F�~1��ȹ0�4n����H�ʿdh@Ϛ&�N�<7��4��cs�g6/��}o�pm�D�a��aԤа��жa����6�4M?l�0�[#0.x�2�4�k�� �+c7�Q%��N�e+ ײIS����f]-c��W�9�	����ƧG{C���^�6�� Cb��R�ޕ�%#T'TĨ��#�!(O�i�7uA��ŷ��p�!�T�!v�7{i�C��|��$E�:�JX 0�̨%�\f%-���>�w��6���uG�)Cj��G�o(�p�)S�1|'�<��}e���받P��o�8�w�͔���_Y���!�l�6o�;-<?�krE�hn�Eg@ցb����1u�~GWVO.ʱ-Z�����G�p���'��7Hmo� �n� ^u>Dc=[��t\�pOͶX9���;F��`��`Q��$Rq�b�ܩ<c���ώּR�p������+���K�m]G��pC+��K�|λ( ���HUs��g�\�Ԗ�2�K��^O�*rȽx/���Gb��贑OewbS��Љ���.�q��/�!�� .@)�o<�V1dD����Cʺy��1�Dce~H�J���Q?G���I�( �҉�
���~�x�-;1ǲD��\̃Ɨ�u�v�J�d��!ɔe�8C"�����7��t׃Xyp��ՠ���ܻZ���s�Oe�Q*��J�M��rj����	�H^�mk� �����cm�MimG�ٷ���Pe$@�,7�\k<���H=��n�G�xw����=�}�c؁ ���u掰��(e20�1�Fg���Y�O�0�N�x"�:7�b�	�	ӣ8�u����E����n^�$-r,k7J�Ѓb��	XD�l@���M���3�)(fl���k6Y9�@*lZ G�{��ZK��d�CfH��<�Mڴ'. �7m8֞_�t8�/���X�C�^L�X/X��������.��1���'b\��E�(������u"�Cy�:��D����.0y0_�1�X��lF-�mNпN$m5����R�6F� ��<�A���c����s����ܜ�H��\�yy��E0�>��*i�_�v��M-���Bk/�z�<=����@�vor�tŐRL� ��M�ԟ�� �6��c/�ٷ#�	l�A<��F�ߊ�~�)*��y�}�Y�[��?׷G�M���N�<.���/UŊ2�Ĩ��F%}��,`P!���%P,|�����
C�UTɋV�*<'̊r�@�8��I���	{YA����o��L���_�p����>i)w��L�/sp'eڲ�J4@c|ZՔ��P���ƅ\���Ќ0�O��r �(�aL��i2R���zj��~��O�v<0�!_�_��y%I���:+����V���̞	p����g�o�և�����N���3��A�B�g8p�2TIL�A�Ї`�"�
k^��E�Ǫj�N���=M��Åyu2�a/&�޿eA��Cb;�<1h�q��2^�e�[󃪥�m޼t�/v���2�)�O�fS��+EKOo����x�5~�L	o��;���������J#����FWF��.��?o���wh(�@7ލlg��詅�8��C�\�*���ۂS�־�\�<*}v��dyw����."��Y��,�ճ����ɫ�ު���N�K�'����g�f���~e�I^H:�ҭ/��s��r��2� ˯�\rA����L�ob�g�%·����ty����(��i�^|���fJ�ٲ�r�-y���^ߖ�%�	�j��
	�e�{��3��t�S��;��q�g������8�����r��
LZ�R)NF^yi{�g�� g��qE�K�s���<K�+$�x�=G�m]޹��qxn���K�u ��U�j���:x
�T���R�t�|�r���w�IFx�wW9[g'����ws�k.��cC�����7�A6e%G�����>A}ra`����D��?�m��O"L�l�L�e0�p+X�ys�ċn�jtX2Xb�7^ǩń��9�{u�ЅZ}�u�!7Ԁ4v����d9A�&20��ݎ]R����E������FF����oδ��Î�v�e��"�z���T)D������|Z�����a{r��iy�8�����Ҳ�K<|ҩF.��q���#�YUW�'�e�)�5?]�:�S}NT~���'�L�,�{`O�[X#�i������	� �T�ؐ��!^͟�J�1���x� �:�� yS�&�Z��҄(e����6ɐ�ti��ᮚ�'����"T[P_���}�bWy�U}�@�O��7�h�'oփ��������� �9�II�_�LQA���������p���Eb�a:x�2o��E$�/��ffƢ�|������8���&�:w\ީ���.���clY�@�ծ$b���=u��!6��1�i����iM�X5t�K&�n�?�,��	�9�N	�����o�bJ�yk/@��$ع��644��@<+��Sh��NV�N$q�#
��\��`u�b�5����k������nh(��G��"�q8,�$��0U�v���<���˂����=��ٱ���e������T��j�Ϯ�/���� ������k�;�|u�-�9�%� �~��(���a�iz��IgRKt�q��d��w��K�	�hmW�<��;�ɼ�x_��a_p�����]�p�ȃ��0T2��z�E��~�t/]��v���X�Ͱ9�ۿ�� )��-���z�¬�ڬVN�Q�~��$�>�=(��A���!�>$o��lOI���h�=�ViTS<(#�)�bǤ������C��K��#7l�"���o�绥(4R�7n7�}�C.!#dӗ�T�m���w&{uP"��;[��t��{Dt�]7�	XR�Gݨ�O����k����2����Z�@D�_���7H���sYm���e�3��ĪL�8�~��eӽ���δ�5�Q"�^n��	Ŕ�qǤ�Ń6�ٞ�s�A�*��x��㈣�=ԍtt�O&���|�o���IQ�����	u������V�bl{��`s�c����R>Q���(J��i�&	�U
�?���T���M_�n�|b�Zo����mE�E 8���#���^�ca�?������h���ܸJX���.�Uz��AR���@�%NOH�H����z���ɧ�o���J��'#�X�9���t�ن�@@�a ���۫����ґԵ��>�$�^E���s5<}��	%��Tt�En�&����_O����QG��JI0?a�"�
-�8{EǏ��~/�ށg*jGGF6��Aţ�/�FQ]�ȣ�B��D�~ �?���-�i�!��N��bZ�+�}y�"�	R��t�|�o�-�f�!0 �{7;'��� ���r&cD�]�a�ԏY:yz�vЇ�%���s�z�&g3
J�yb���3l�^���?�mcYE�Ǐyԡ&�m�W��d��"j]��4H�S��7"�����nL���,�ꩉE@����)�_�W�V�fU�@KN/�J���]�Ť�:ϒ8?�	>��:�"%��č �����0U
STg��lP��*����'y�Q� �%BG��DXb�I��s���e�
2e��I���Py��g����l���8��4��}d�yMnr�!|qWH�"�BV`0�k���X'��l��ڄ�
���?�Rq��-���;3|���'����j�qg�w2rr�7<�jK*�o��tI �ذ.Huv��{�P��9}����~������Y���e�A�������,��V�4{�e�F*�I5�2�!��k��5Ö���%:�T��≻�����Ci���T�<��L��WlSK�&w��a@c��*�ܕi��3���
/s�LM���q�����X�H��!ᗔ|W�f�uxT�:�\�=�����M���ӽ�@vcc�_V�>rr]��YJΛ�qߠ����VN
Q��̯��΀�p��&�m�;�F*"|}h�{��.�;<�F�R}�� ֮�*B��ODJV`�"B1��<�"2�7�K�ĞoBw�ȅ� ��I�uOs�i�y>Kw/{�5�(̜��C���G3�,[��?�T*����V)�u<S��ߨ>|�㥄n��v�`~���$������; q�ξu*n���nD�W���X���&�HS̳����'���8E���	-��?a�{Q�-o2���j���ĄR�m.� �@�a$�2b���rf��/I��� vԤ�$s�}x1P!(��ߵ��=�z@���U�)6�i��J��Rޝ�[R/������[�h�5B_eqΓ^�S"C�tQg�6���O�������t�[O�#ZG�۔*NÅN�Y{���L]m�E�n����k��vBpٌ�c�����tbչ�%Mg.�:�^o�Ӟة�^��˓F!��p�f�:���J���jWV45��U�]s)e���?����ŀ�@����09���NTq��ML���Vl��K��:��ir�Њ-��Gq5����E�L*Y�b/�ť���d�n�+~��A$&�����rÞ
�7ok����}!G>[/(C�z�f�b��aK4��f,�v��`�!�T����8P[q���XO�`_��x���ڏdi��-\�οgK���;OKQ�7k*�ǝg'T�Dȇ�N� x��H���^D�T�"��5Mw}QG���UV>��[M�EE���'�Q=�୾����F�߁u�� ��O�lpbҫWj e ��<��*!�*r�3s�XB�D&e�J&�1���[�!���{���MO�&�:S�j�s��=���#Q޸�gS^sÎ���լ�Lx����d=m|%��>|��~OP�E��y�<:�ovҜ�Q��K��E2����dZ�(����h�C<WP���%qbgr����3���嶀S	j ;rx!�ka�]�LDo^�T_wq�"iG1AK<:�0�����Ez�v�]�'��H�_��=����g���������0�Y�X�)����g8Rp�[���(�-���+��MZz��������k���R��,��OKh+�_�)���-�u��M���n�MB��Lr8'oL�j���pN\�:�C�v��.���yN��&+-}���ؚ	��?'��.�KF]��yz4ZfvO�b_4��V�L��he�U����.���R�I8_p�x�Ls��Jzj6.JMl/�T����h�������o���$��rRX�'j)D ����^�R`�7.�d�E}"@G�7���6�j��f�xRz���{Q����ζx� |��̠�`̿�%�GGGЬ����Z����m��J�T�c�,�'Lq�YU9�n�Z2߹�9�ݗǾ��ܰ��՛�D;�<ţ�?��YH쿋W�sc`^+��>z,�#?C�h��[6���	�đB���[p9z��%X�F�p6S�88�Dɷ@�a{�z/v��ҧ�e�B��D2q_�I�Qk2fį�1�t���ǻ���yP'�̟"S��V�Z�_�����s&�@�mN�O6Li=�v��J��dx�?W!���mQ��^����Iȉ\ȸځ����T�e|�"	ӣ.2HUg�����J|m�`>�����a#���7�=�kpAu����f��@MmL�Ŋ�76J�t�"�[Ht)DZ����bolX�{$�$r��w�^ļ���Z�&�^�[wOS{9�)��.��8v?�b��~i&��C�I#��}�/�p���}�`f�])��:E���.'��EY��3�H3��YG��k���կ���5����4s���0��Y�.܊�>[��d����yR�����%���%��*4��9�4%�� ����%�Q$��l1Q��D�X&�xw�7<�-Y��# �]\�؍Bc�&��z���å^1��7κ��2�(@��� %��i=����&��NV>�*cLIZ^B/Jm�ȁ�N2u�W�r�ڹGɜ%��񭉱��mh����3���&��
�,�J��ڀ���@Mo#� I�?�l�i��c���ƪ5I��t�Rɢ��~&���6���2N$�0,z=W"?}U��lɮ0Xj�������*�4X�) ���/\!��œ�[C�u�a��֠�`�ٔ� �3�M�q���)$��<=�q��ӂU�Ή
�ݙ��_o��HJ�^8�r�s4G[e��|��$)��r�b�%��փ<���O��_��Ϩe
��@�vA-u�W����e�ek��6����&�rvW�!o�?�X7�-�a^Q Z���cs�^�-�@<[�����_����_���	�d�9�`��	�2���^5\��0��a7���وe%������Z'���-����>�px#my�3����gv��\DC�gg���a'̚���ȵa�ui��JL��]yc|��'4�R�$IV�/S�Ԉ7o�h~`!�čƱ�R��$&'ǌO�'��٥������&��l�7|^��Yo7��|�̎J�{��7�R��7�n� �k��&��*�m�ru�ð�D�\F$d*A^��k+��܇-n3ͧ������Λ�1$a� 䴖���޷7 !�+�J�}A-��^����>���-2�w�6�~�}�x&�ݫ�ue��{&�ȃWWm*�����Z�s-ģ�ĬDc6�ĉv�w��ҥ�+ԫ�?{'e�X��=��U:5���dS������&Jsi����E�!�rQ�f�	�x��W�WJRƬ��pG,���Ѡ��Yp[D�+�i�%���WG��-�3���%�v��҅�樁�Js��,< �Y�}��)m�l�9ʼ�0ʠ]��q_N׽�d=*����H���_fS�|ʔn^J����U��xy�~i��b��\��|Uk�n�!St��-��C�N��cu�@�ͯ,r�LE��1��CKjY�Ѫ�䟈��9���j9b�_���2�r&�{���aF��c2�k����.��3���5�F�2�T�/R���#���M�G���S�6^7��45M�Q��.�Foe]�Ťlg�1:�py�\�zݮ���T5X�%~h�ٳ	o��atk<ʆ��z��n�/�2�­�Q���oۮ͑:g�G)�h�.b���^?@�8�Ӭ�)f]��5���E����L���j+rU!P'Gd;���ޕ#8�9rȏ��� �����f�R�S,w���q��-v�NZZʔ� z���#�^B#��7�"�rX���o%T�d� 4�p�`�[|w�R]���1*N�n������M�w���Fl�����9SR��|TT��S8H�� (&y��6��'%��0�I��!���-�,�D%����� �X��q����5�s�j*I��_U�@<~���~t�f�q+�WH����ĵ)�C����{Y[]�t� �ק�B��C;#+�ʱ񹇯ί��E�g��/R�`z��eq��m�L3K���A�?O|�O�l�d���(�Mf����t[@��C�W����Y�S���<��毼b�M��p4\�� s����d�2��ԡj��sB�źG�K1�c�u~����`/�I�ӕ	�eO �r����^�8��7��F!�px�'#9����z�例�lBw������I�����tE��R!��f ĘbzU�r�+@y�v�c�>S'���HHryGP1xyY��<�?��n��R�Ҏ�?���v��f�?��=��<��:�s��T����u���f�Òf���3�3,h�F]Ք���p�^_����M�CJ��/=^����qڱ����w)������|�:t�|��������4R�5���(���u&>�����`�P�	-P`�����9!N��oq%A}|�]�}�|�ՠ*G����@�\jR�h����6�b�1�Ԓ�E���~�dcU�_�aIn>&��>����(��+�b�a�Qq)P�x_R;�F+��)��)F_ 1ۋ H܍)e��>.6�/�}�Q�Q��1�-:{�@�	WeE}����y�j�b�t�g�!#� ����&�. c�c_�}02`z�nzC�H�n�"KY�7�ka���Rm3�g	��<��hL�U��u�A�g_�kՊ�>�4>�yg1@��qGT�9RZy���Iy '俺n�>_�l�pJ(^���'��Kya��_zڮ��G[���F��^K?Bh*Ptd����{���h*�Id�T\��
��ѳ��� ����n��2X�i�\g���hC�Fy�y�a����Kն������՞��*��!}��NJ��_�ܲa�32��NM/�5dx�u�	k V*����4,���A!r�1��N����~����	�����l��}e�Z�X��cإ*Z�+;�Ut��u�AUgo52W�6��_p���/�_&��s�a�B�x"�h�s�Ȣ���>Of��"�ͱ���ց��A��	"�p��Nnv\1L饩���|��n/�h�Qo�tHy��1��w���P	.�ո�z#n.��e7Z��;�@X02�r���;����\�WO֢� @��(�ƽ� i�d�;%�� Z��c���r�������,���;w�<O����:����0��ފ�R6�����{&S:�=��<��F���J��,�U<dv	S��ձ����~�k��҅Y��(��UE��j܀���?cI���d�zpj�l�y��0��N�E��g�ryI,�YZ2�1��!��=8��N�7�tuO�0߃��lBPhjy0��5�����x�J��_�lȲ+��R��)ɊIU�|�5�r[�/��	*��,^�[J��uD<a]���u/ �X�l}������y������R���73�'�R�/LPRewXOӫ�����8,I���ѩ������Y�xL*�Ԡȍ��C�~mO��N�sc��FRUp�A����V�8��u��~k��/})�t.�9��j���k������S�vr+s�Xe%�l���Ha���WO{�rI{\�ZB0��� <���y��rE ���|~�D��/�LÃ,\^��`U2Z+��1��0o<��yZ�Y�~e�y
�Hh��}��Y-
/�پ�	��m�g��{K!?��8��'�g*x3VR�6��j0�mӿ��I�4�Ǥ���$�l\I�Y�������1�@�m�^2I�END�L���i�lƭH�$$nh�n�BI^FR>�"v�ɰ�G7��gC��cg�2bzO�:K��V&�����Yo�����n��8�T�4{�Ꮶ�8 !�,ڊJ{i����@�<5r`�eH�&ԼM�.S�:�s��;��Wr3�`�gu ��s��o'��x��.�_ni?����v�;+�i��۱�<�V�]N78˸��q�d�I�� #t�E&�rm� a���b��9ϔϔ�����[����(��G�UW��RC�;�b	L(�G\�M��[���e���i��v��Bя�̥�ȻH#�1I�ڮl)`Z��
�H��iǔ�	�6�B�Uf�mp	�H��