��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-kc�wL;Ɓ{o�M��	1`��.<�8{d&L�Vi�,�ڠ+�\L�������nv�y��w$Q��HO�_�1�5
�Nt���7��?J�x�*NW�dk[�Cf��6M���M�oW<i�("�F�<ߌ^*�Y.���{o2z���/����Y� /��#��D�:�l�=c*�G����.�-�Ѐ~����zk[�~�l���#���U�z 8�:I!}B�B=����ui]��Q�à�r9���/?��|��ǺK�뷹ͼ�5�"���ޑ���=oAV�5�2,*[�GǟY/�r�
^�7��o���Y�	����j�
O%��.���Eϥ�SJђc%9�����16؎���f�ܯ_������pk0�ܾ�����$<����J@kY���0�R�F�Ci N�1R��/�[�,�B�����y�
�s{��_�^(�-�!L5s��D�Bw�ɪ�}�e���jR��}�<xJ�-5s��V��O���/��������q�Ay뫠M�(';ui��W�n��U�1FP5W����;��n��hFV�\,�e��dP?�1!�m�I�5��;c\H���r>�c[�� ys�v��&�
�֪�qR�z%�.�&v���I�T��
1����z�A;����7���},鐣����w��B�ݷ^?��2B���mdH�yK����d�_�k��	ς�`-Mj7H���q��~�-Hj����[B�=/�8�K$ ����Q�f��ҫ)7�SWy�J���� �L�^9y|�.i9ky1���ˁ���D E;���&��	P������#��S^^:�A�Η�|C �f�^����8����<���@�s�t`�50��Y�q��%��{�;���G���6�V��7(�"��g$���,
|��Z!*�Ȅ!����"�L轚�'�H���^���a���u�'�	��)%g�����Qn��H�\7C��S���p�Sv�5k-��(-�qo�\,*��#1�ަ.������PK�u'f1끲㶋�:R�2�D��T�/my*�-E�H�k����������X%�|u��<� )Y��m��-N�pd�\^�k�Ê�CV��'�&H=J��_�����N����}�ĂN�+������"�F��td�G����߬����B�S�*[���	��gS�Y/)ȕx�)t�V�D8P���_�a^g����0��f��̘��j��;��	��\v3jm�2g��`ǻ
�e9��R��g���-�S�����Q�Aշ`?z�4� I�h�R�+�����G*�y �I#��kF�:��9���+GEo̮�N�'�w�3jж5
�Ԍ��-�v+���{6��u�2�~Ƞ�Mo{��e��U�mkH�f�M��l�M��ە��l���b&NT&�J$�J*�b����f��;>��s�/�
nV�Y-Q�*>�
�'���>�f������:<0%�.X����&'����T�PJ�Ԣ�M�W5e��9��Ȼ�2jW�;��:��~���F���Gܸ����H�.B�h"ș�wP ��D�A��7���}�Y��-��{֠�3�34E���a�.co8i������=�mIR�K]��cUz�ķ�e;�XL	�K2j�\��]��/:up����� ���A�	'�x��f���ZqY-�R ��9MX�\��&��Ҵ�ޥ&uPFWO��:�\�UEF2�B �\5b
��(f�x Rxs����V�\���E�s'���Z�y���y��Br7��Tg6�fХ@ۅ4a�S|ɀK1�� ��.[t��x��K
�X�6�A�	X4�KO�3��D�?N�����z߈�ן1<| ���o[&A*��=�����b�#�j�D��C(�,|�T�*k/L�-N�dQ����Rn�ہ������R���S�5��Q�Gɶ~��O�;ǀ�H2�d��k�.@h�4�Ú����~��m�/�X�Xmt�$չ�R�-���^��׀��wO��,��z6�o�Q��|�J���O;W�,��hT<�m
���Eb1m�$��2iSj�ZA�"�r^Uf���q���$�_�,����C������@�zz 2�%C<`ɀ���!n�$@�_+#�^�<��0�#߲9���j^4ߠ-.�S&��YB)�ww�(�*��s���{��n6����2���z���a��t�u���^*�{|����=�����!�����[&]	�ЭO-6,���{d�f8�9+m*P�5<d��}�<ݨ�+����F*F	�;G
!(v�V�����i9���RIy�Y�	��%�w� �ٵȐ�)�qf#T�b�Ӧ��1ΠC�tWCd��tLr,����6,Wz2;�I�V��Ǆy��0�Ig�3���)�9FȐB��d�<�"�O�X�*K��@���*7X6����ڈ����E7��!gl���BM�(�:`"��`�?������CP]]9��x�j�)x�S���ޛ>��{��-�_�y��|/�t*���}�cQ��䷎�륕vB�`p�}o"�+Hf�8�="��B�ra�j+�5b��'���@<�G�9D����ȃA�-�ˁ���6��Y�@v���yYm#�~2�����%>mX��c �~�
s�@g\t3�ַ��`�p�c�q*�?����mb^^%mpE�Gg���Ӫ��3��!v�IMII'N7Yc�m��d�x@�}�����ӗn��uܪ���+2���@qd!��1'xT���
f���O?��Zѹ�������?
30󀖔y�5s��_���{�A ��Aߛ��,�l�6`}
V����ud��/��ڷ�w6<<R�-�j�>�z��AK[�ۃ��PzN�}˩���vP2����ʣW��>�R�|�t�.5ng��E����0���W�����g�U�f7h	�����r�:d6\�/��=�z����7{R�h�6�N�vPD��S�T턎vT���I~)S��sZ���g	�Dq�&����]�H�o'�g$�u�	����O)�Rm� ��*e�O4o��d����ӹT��S�=����Vb ��=a`L�z����4��L��Ɗ)q+�G��l/�.�Xe���mDAI#�����~� ��z�~�i��$8�A�IG���8LZIшK��zyY�)i�j���7���GEj�ǻ(=�5��Ĥ���T-��A�1��R�!�@oq���k�S�ۑX�,'��/2�z{�2�[S�4��Zb}������$�xRux�o�Y���HnV��6�rKv����3�nPx�`��DDq-
?��zt����ҐL�-��\񏏏
��"�5҂*˪��1���e݉@rC��O��JEG�y*� ��0�쿌/�T}�\i2(��	���JmA	�Njb�cΩ��O�8�@����#u)k{����$����Z�>�Lz�ci;��^���-�<`�*^E)d�n$(��jI.#�nOA�q�N���0��{,CE�]ډ�x8��E7"ͣ^�Q�H&k���`�Ww@X��ѰJ|����6�07�	ը�7d�J!�����9KW������ɀJ��/�V6��9��\U�F��v�00����d��']]T�֧�u[��i���~i���o�f���Pq�Q�6�F�t ��]�e�k��n��qCE�f;�SmJ�qU�a+�0sX�㼒UÑb�CO���1��C#4�f��HqSX�'�PW���� �!���6w� XLvM�?մ����CZ��X�Y���
�ڇ�8�
%�/�Ym8Uѳ@ٵ��֎�k���ҏ8���MFQf��g�o���o�T�=��]��J�1?��X4�c���V"{d��	 `'�^r���S��gLG�%�%�����17�+���4!xr��TeW�Py�^t�hQ���[�
u)����L��J���n'U��=��s�9� e��F͓�,���h���H�� )�%P��q���4ZF<�9��ݸ��2�����y�8�c#�/G<��>"�q�]�R[�d����ѹ�~C3C���}��&�#س�Zbe ��qw�y�ywzW��S����۹�-)��o>e�6qwL�C�K��P�D�˅�X���")����-D"ɗ������jA�BW=��[Z��ms�ѻ���WQ٘�w��o�'=��T�;^������'���gN�H��������!��܍b��P��y��R{C� 2�z�>Z+��P٢�kI��!i���b��3��ɾ�#%��v�é�y�ƽ�H��S�,�/�YQ�� g����k�̙ΠJ��z�j��yE�,c�wn�UT��!%`e��-�A�������up�5�궟�jS�1�0�6��u��5�
��Q_�s�����fm�����2���lZ��ܷI����ga�N2�咃�"����w!�St7�5�l^ Йi1]�^�ս�qu|~�rn5��iY5�Մ
H�id���s(�!taM��"j�Hge�_*Oz�,%�ũ�C<A	���l	��r<�%�:�#O��쨽n�)���7w�:���w�2���i*�.���̨w�%��i�TK��J��=��0{@���6V���1��iЮ��@t �C��PUL�ľ�2i��C�Ԩࡌ����?M�Ȓ���ʓ^AB���)Yd�Jg�l�҅�2e5�_/ڤ�ņ>��M;襾�Nӊ�N��!�:�7��4
]�$�XP�Ƨ��]@j|������5�d����O#M*7�_�x�i�;X���ݖ�)�Jֵ� OP{hcm��X����e�{$�m������Z�lvr���*֢xĚ���<�Ð���9�z�-�r�J�ᥳ>(�/�� � Z� I_�tZ#3K.8�Π\��޲]�m��.<��;�8[�=�T����f���e�QO&���fCU�t'm�%���^��a��~���gJ��.�R6��/r�`x6�prux�¾�l�XL`�z!�^۾�-�7Z��r�؎Gb0�8ިp%��D��t�_*L�6�m1�Hi n"�\�-��H�� g���&G';��8�B�*�
����p��q�����tFG[�^s��쌠3�>�e>E[�m*���S A��M��Rh�)qФ��a� �p�T��l�N�$���9��t2sy"��+B?�^r�o�<�8�+Q��]��W�	��afa`��!fHF���c!JDa�m}ʁ/�� ��5 .�@v�.D�H>'�&�� W�K[�<���?F�KC�k�>ӥ�Ȧ�F>�A��5�4m�b�K�Wo�Qv;h��1�g�MZz��U)��o�,���?
1_7XB*��˪�ѧ`�'d�67>׬!f�4A%D�8!��_-�}���#�q��BLh�7ļ\i�R,��A{��{տg��|�D��}�EC?y��֙@�Y<��G�!}���h]��V���֝��C�j���n��lE1�K%��f�kEp�� ����jv=Ƀ�}�2�]��
�P����?WT�& �2"�G�/��� �#i@�|��\c�1*d���F�ج��=d���<M(��Zkt8�Ҽa�&�(_���Sp<�:��{�E�X	뚐�'�`��`���w)骇���^�9{��p��M�"�^,�0Y��ı]%�/�g����0J}�{���
����<��Z�;Gz�ȚkpZv\���f�2/4#iwmW�+J<�2/��ܔ%���w����H��?�^g���[����i5�k�m�r)s�*��ա�f�ي\����6�۞
B�A��/m�{C6���\�ՀS��;�mX4�゙.tkRʅuFe�R�/#�j��OR�E��i�P�K��c�sr�$Ntr����y�J2�ko�n�U���	�sT�d��؂�eM!�=��9��[��NS���h����s�Yȧ�F�p����TB�nd��������eB��i�/-��b� 3fa���ͤ���p �s��:DA�d���4Is�����hWf���A{�;6��F��T`��F|�:g��/?6I'0���tW����>V�"�U=��R=o6���R	��RU��
0��#�_ BD���D5\� ��^0Qϥ�ܐi��B��bN�"�Fo��?ů��w�J@8A��g�hs]ȇz�6#�X[��0����<0�g8�-Uz���v���q�9m��I/Ak¹I6b�*�bgRY��_����0�Ud�ϴv���8�"	_{cU8?�~O8h�ؠ�^��9�W�cRnq�)#c��مSR�Jv�&���Nzs���|H�k��=L6{,�9^�F�;k�V;�Fo��z�U���&��f�3+�W���D4��Ѕ:���cZ���	��!���?�B;p���r�D��
49`�fY���S��(��d;J��	Df&���9F�����Q�*��+�t����x��*���V�1�D$�4���wT��h�cO��G��]fb5%��1����brba�D�y����<�����
L��
���jڈ�$��fY»�m0���X�,��i�׶#s%+q�Tb�����+��εd�>:<k�j�̚��g����ʧ���I-��2�ܾ_��V��-ŸWBe����2�=>���N���琗�����"���M�a����a8{�E@V��!��Q�Q��oN}������`�_|O$�E`�k:�G�n*`���F!]<o;鍕�v���`oP���Rk�A_\���к����4�w钓AeL;�>d��)�����9����E����y'_s�Mz4��^&��xH3��j����g�$̳a�xɺ2�;z!��\������:U����3���$����=8��`pOE�ެW�С������&'y�?��� WH�	�u'W14���-F(d5��d�T�ѢG�i���_R��d5�̌�C�gg��(��Ǹ�~��6�?`!�Vt8��'�*��b �]�j�SYbQ�o W�]�=L@�����n�f��KOme��^��f����璣R������t��.�L��?����� �����U���L�PF;O8��م5nF��@�8��4����E�Rv��~y)��^Y���)#¬�-}D���E<��@tީ��.�|�pе��;t�S�~�
D3�sj'-��N���b���e%0v��qK8�fz띝�C2��Uk��ka?�7�G�����zt6:�%rfInHɼ�nJ,F �F���Li��$g1��YB[Y��KIR����n'0^8#֊�M.�zxyq�nj�����u�V�����X�>�F>��bg�+�fť��x�y�c!�]q>u���*j3?k�Z��R��Q�qn�st!אyhl]�j�����T��
j��H���M��}�`2��<Vժ~A�Y@R׾�$,f5��;���%�^��d�9����� �^�'���(�v@~7�YrY�@w��TC4��Btc:˙b���W���6Lal����!�����y�'5�y3i�q�����Ǐh$Y^$���(�^��a�lW��0��t9h%_�M�,i�@]2�p��� ���y�w�I?�Lᘧb¦a�H�M�Uv���4����4�v/V!a�o�|�.�b�dt�ƶ�=��<����9
��1M�C�c��+�V���=����ѿ@}�.�Ɍ�d�󌜣�n�%B�k:�+O���{��PV�̹Q�DiZr"���7�X�p�h�R��?�c��Wk��NT�����^]d�2k��,�P4��X�+���H?a� +L҆uɖ4��J��T<E7��o�@��M,x�/3�ǂ�d���k"�<��Lt(�fBp�yg�'A<�a8�zR�ޚ��U�!MM�c��,{x�E�dȀcں�Rʴ�ps8����+��,Т�|B�{S: ?�R�����$��=����^]��4���ɹ�-������+��[����yXo�!��ہ��/"U��|r�L���xu�6^��n]�f]�TS�.�3��u�����Eq�4�p��6�dU���!��<`�ڲpa��_���LÆd����p���mBA�����k��r�7l����^�!M���XI�>ֽ��g��9f��1�M`H4��3#fu�s��D�g	s2 %��#�i���U�����ua�V}��Q�;�]�H�w��WxP�|E���J=��0v�71�pkҲ��O(:��T����0w#�8c1�u��x� �W��G3��p8� �$"m����b�-�g�a-�^/��C7{]c���/֫6
���C=�h�Q`��(��r�8���T�+PL�Ma��Y�5g��C�c�9��l`R���k��?���*�;|�	��}����P�F�ue�<b$�#�l����R5�T�r���(�2)��O�.]�nkVh�j)�!����0@���+dtߡ��7Nw��U76w�z�v��|�L~Hl�I����Δu���!��_r��ra[��&'Cڂ�5�i��9��eK����K����j��4�;��2�CG�U�I�>�^�$2�195Y;�m��@�Y�4Ŷϐj<&,�gr�)���#�o������rZ_�>����
ڰmJ$���Զ�D>W���:���_Ks-,���{� `t��g�EҎVjD�.w�������A�Z�kB��=����ȏ�D�?P�,%�:5���)YH��^�9f!2�?�h��G��^<�o�]��=��*���?gՌ(c,�Ih�d��5#� z4#���j����<�n ����yƋ�H�r��qJ�A���&#� �M���_�Xy#�zr쌌���Y��N�+�\�zo͆c^�$dLl�}�Y_y��Z��<e����z���iͥ�t(��=]��y�i�р�ܤZ�,�k�[$�uŌ冹9A��c��V�_Z��K�EC-�*yΡq�lX�8�����g�3P
����s��0��f�:1��Y	����A��v!����w.���:��5'_�:�1._��j�1v$��ŋ�2�����؜yx�ݷH84�䠶�<L��],����r�ˋ�*�_��툻ʈe�48*�7��@��nQy)���~_���||�4�[3''W����ɞH8�C�
%3����h�R��&8$,b@��n�	V	�j�6|�"jK���H�5�|}�q,Qwu�x	Dm���`n��߄`��B�����p�RK[���.|{Z��Q"��Pe�Y��{��D�QU����DK���[dZ`���98ے�ѴC$������ӻ��~AN&��i����J�9\�Z�v�y�ɫ�Z:g"p�隐���4
?mBo����s2���(�Ϗ�l3\JT?���dT ɺ�L����@[���\�����q[jul��q]���/$��6yQ$�H�ov��f!�3���O*����>��4ϱ�S>�e����.�^%va��V��~Qc��E�Drõ}2Z��'	����C=���&�8���0�C��N��&�%�Ld)�<c�n'�cxhB/
T�ݔ���ICGqKY*�g�]�Z�2�a�H�$wo���.��R�tɽێr���aJ8�7:��c��*�b��t�$��]/^�?=G��0=-�3���	ٓ\�AE�+��`�o�7&'������VF�`I�(�(�F�3R���X��LJ���ߛ+�tJA<p�W��wH�Z=��/[�)�HT"-kS��1�=�뛞���xG�9� ��Q^����p��ap:��lawv=�;��Xь�� ;Nz���ݻHr�����k��U�Om�}�8UG��-2�n2�O�O�,��d��8��~�*���¨���	�A�w��Z�_� Jy�١��1pXu��j�m7�> �ɰ��n�d)y'�D);Tp�\������0�(H";��t�K�m}�+��6f�nZ&�N��
Ed+Hh��V���H�S~{����d�P�7���>���"n�w�bI�Tm�YsE�ڠߧ?���ƮC�і��?����)N��8�~K+�C�Q8@�������7��g�2�ѥ����p*J�pxG�?����G`���Iy+�3oIK���p\�J{���d[_^'�AnI��j���ᡝ�%�O[�2n��d�m�^�T�$y�ۼ�������ˋ�M�+�6 TdPn�r���=;lN���e�����c%ޱ�9d�؝M1�.*�g�J�MI�>=���T�O�/i�iE\���=^��9f����)�D
O�E���2g6�����N1�t���gn�T�:���vAM����
�B�H��T�Xl�J�T�Qt���k�L�z0C�-�D<���ZaIl%t=|��A�Jlu�FiUV�`5�;bUX؊pՠ/��"=�EA=j���=����~�X�y�ɞHmx�/���"x�y��7���f;�������s-���Dku h���/W�q�5�H�b�a{{a#e���~\��j�VdH�1uŋ�<�?'��AD��)��Ac��oz`����Sn3q���F�A�e8�Şq�p,�f?�Q�*��!~�r�f�����޽��ez�#�a���:��7�Q[~mkEщ:J�������4�����{�vwS�w����1U������-�FPU`����J#� �Q���j3.���\��̏���f�w��OgV�4����2[=����2\+BiƜ��"���6�Zx}�V���D�l	�M
��f	�Od�y�iV�`\Za}C������p��6\�x�h ���2���z̦��&}��M}*�s��	��&�{�X�@�H����VŊ� є�D�d!w��5��˹���=c�[J�i,���Ll�.���N��Xh�SeL���dƒqk2����UZ���U�U%:1��C�������Ɛ��x�]XcI��˿���߯
�M��7���!igPbg@�����:����e�x|0�������K3d�I��A���(ASP¸�<Nl�	���)�T����n��A�U�G���'Tl#;MT��tjqh����5@#7�YQ�'�v�}Ǥ������	 Dr�ֻ�bU�;�vG����R\&�X�l׫��`R,�ǈ��悂^�J����$J��"T��R?a֒�v�(�̼���@�fSϷin���*8�f�f�솎S�R��M�vFg�Rj@���(���m�c4z9��"�5��م# s�۠�4�Em�4����{��	��mn-���n��^�(,�����0����:ԯ��P���,��t���V�-|!�;�F���Ǐ��4����^g�mm�!���k=�N>�������T9\��N'��>��F�'~�ͻX�Zu&���廰
>��=JS<���)��
ג|0�@��0��S�./��&Z@S�e�#�7�'�-z�!Fh���\��=�-����8d�1+΍��nѻ�>���p��ٍ.+ѳ$����P+�lW#�����HkO���p��,�`�iO>����������U~S�:�+NĮt���'/^%��X{hN� ��Q�N��f�y�����׵A����h�jUv�W�����)	 A!b���pFi}a�Cy:aW��Yߔ]*.�5ɩ��B��s[[7���3p%����w��b:����I��i»S;���_��S��Q�o'�@����.[��l5B9�oa�:�X4A1Ԧ������FF۳c
�[ �V��,��ɒe���dƆ��}��+���gJ�i�1�$Y���nࢤ��^������0�t"�o1>˟Dhw��A.�9~,j����z)��)��{�`��u/F��٢�1 ,�� �CBr!�yR���Z�j.�C�E����9�*�ڍ���ߖ��4�(v���m���*���9��Ab{x����* ͞���� �Zи��9̯�\��v�=���[<���!/Q_n~�V�Т���O
����w�ș<g����*�7�r�N�=u4*-Z�Y����k	��e�/��X���S�G�*~S�����ŋZ_J͓1p�3a,>���)�j\]!�P�:ǚ����|^��f��EH�9-�FPz-6�^S�zH��Z���_�R�& ��܉�ať��d�6ɹ���C� Y�h���~@��Teϖ��t���
�It���ZBe /y ���F��b7�!|�
��@ fm�ڈ�/MA�4-i�	o5Bm����T?�Y�o�&�M>�G
��әZ�Cщ�ꅉ6b���k�8�܁$�V���"�M��y�"d�C�����ԏ��Q��`#�����E��K�W%�d6!��g�h"w�����3b�7B�vOw�9����E��ud�����x�>����gu�Ps����e^o�+�I'�]e0C� G�����8Tw�{����M�]i�Y9�NѪS�fg=��=��������+׼�w�c
QR�/������I�,���u#��뇳�FF�ӿ��]�Ϳ��!�?���pyc��p+�5�9���Q���m2~F9�P�*D�y)���%�4���je����vte�as�i�~|o��+հ�C��	�͜E�J���=23�:i��/:�u$aul��z�Y�Du������
^0�f+ ����g�I�ϛr��UL����6�K�������cwa�����̠^n^٨�����"���-�x@s�Wg�ˆN�2�
�"J��)�g[?��\0҂i�U4����@��۷���T��������d����_�MdY՝�����7��U�7�*�$�"x�P���<��	��y�i|U�<�������Q���Jޫlrw'ᑰ�PL�n�0#�ȱy'�@��5�S�R� J�{���ѯ&_M���1��I8�tC��1�H<x��E��[�g6I�J���w+LJM���NO�1�@E�g&�L}�r��3�~�� /x.�H&>���y���堦�iO�O��߁�J<��SX����r#���ȿlV�"mU!����Q�6���bkM�tE_g��-%gK=�p[2�n����[d���һ��ƃa1���R�u��)�"&�N�w,�!���]?q���]$;`��,�����P�ܥDK;�/��n!�J>N\���d�R���w������.����"��:a�h�h��ʂ����Ƙ�b%�h�8�1q��]}����;�-����0�7��+ X_�[�ݗ�@u9,
�(7���C�F�"õR�'H���A|��å�em�ks�߽@?ɺ������K�(���O�1��5� ĳF|9U]�.&�B!G7��9Qo���~��Z��a��x11J2�M@��WC��:���h���'�y��l�Tc����"���fkK�Sn�+å=vj�b�1+a.A��� m�u��%<����z��c�p� Ǉ�	w�UQٌ�o�"F�+�F|����[j�� e�~����>�*~Mk����{��
��j}�x��'�h��ӊ}���]${�Q�S�"���dxZ����[9~������m��#o�&<���Ws0L�)��|<*lqp�ͪ�g�}�Q�X!���LL���|�����W>��Hi6I�YKT.F<j�Vq/N�h�?V�ؤ�m�wL�)�6 y쵶ſ�ļ�8�O��������R
��pAx8q�S���6��狹"0l���������bE��8�͔�8ځ���"o��@��J}=�3���W�	�:_����}�����_����q|�vɾ�D����b�T�VI�z�h���&�r���p�a�5���%���;MK_`��!T��˲�b�5��0�a�*]�-�?(��:/0f��Mԯ�����b2��H��@'�a�:�kKa��^�~�>;b�	Q2��ei����F��q3�허~<@��6��s�z�1{�6��4��B)���x7\�NL�����x9(oI6���]C��j��%u�����fV$��!���ŅP'�ʋ^�fh�9*Y	2\��f�̣�<��("�4���	�X��O�y�X�	Ri� ��/�v� ��"�U��J�b��_��I���~nI���B}����FW�Z�[�����Fyh��!;�9���c����{�}
�����:e�K��Q�F.OT[���:���[*��Tscw#s#:p�r�`@lq��G� �m7��Z�2+�@V;��~6n#n���n#��x�?6[�aE]@��D�d��i��`e/ ����A9��e���lރz8���u�� Z䔇h�M~~�\q�n��D<0�u�1��L�88�E�)
��U��L�֢��T�q�!WhR�*0A�E_p�0�4�)�\��8�{-4�Ֆ[#��&����Wo��1Wav6��/���G���e���L(H/��\N�ʽY��Y,��3c��E�{PMy��Cl���V	$�xE+D���mVTsn)}������.��9���aN��%��u��XʥךAT�2î�&+�!es�9K|�z�e�n��4Ò��n�`�@K�P�
Y6h��m5K�i�#R�ű�|�LMu��3_M�5�M�HxpF�E"��4��N���ܹ�j�uP�V�j�Y�Cώ�߽������fWj�a'q�u��:q�n�ӹZz�'�iX^:W�{(�U@x�+��W�����{�������>u���R�Y�2o �Н�e��$^z5P� ��o#o����-H&تk�\��m���)����$���@��c;�8j�Ku?u��uI�xz�S������',�D�G��o��:w���໚<2skTx��_i\��;�	�vq���s�脎@�(��9=���vh�~�*qX���K�нRYE��T��e��`��ؘ�S�;l��%ja�M�j��N�0�����2H��w�p}'����Xbc�(.|��ƺ��6���DL=�l���
I�T��<�[�1z��#)�Z�mk6,J�	CCc����7oP��v��G���ui�R�hy���a��>#���� yjBem���Z
	P9K�����'͝�fq$��p�E�x�/1Nn�j����m��ϙۡ@��>��mW�WG*n����&�Q�o3ȣ �a~4|
�.-����d�]�D%!����1���Wb�Z�O��%C)�=���V�>�1�z��p�==zX�� :�36/�6�F@xxaKЎ��O�K�X�fIl��"R����N�6-�	�J��F��Ua�^���WJ�˶q&g���A; �F+W*������^�-����Wō���Xo�K,���MT��.qg�?�=Y���Ӥ��2[�-�����tp�^���;0�/˄�f����c�F��:_1=I{r��q�0?�u�S�%�~˅)O}Iz#����hNl4�M�ʂP�|XW��t���)ӟC �a���sB,�x�!9X�*=yt�a�휘�ӟ>4�&]k�lȌwT��}fxb��U\L/٦.'w�2�E[=D��p fV�;��}t��oIu��G!đ�T��>��[��#����ݽ�s���ƒᕶ���^���j�q�](��A���G��"տ����I�>d��'��O���]���u�(�|c��{\��z��V�^�j��ˬ�X���` �(�C�q0I�#�q(��˂���~��W^4�~L�F%�cN��P�r�W��K����n���\�0'! �n�:��z�%ܭ��}���V��t�K�(Ls��m��)��L�W��
�5�or�;�[tzY���w�w�0��j�cHL'�L7؏Z�� =�����_�*�L�xO�RC�z���CX_I`S<�NE}p� Ɏ[S
L/ɰ�2P���-m;��CH�V[(j0X���]U*�{���^~w��L[�-��m�0_x���=����k7�wV3���v�P�����tG���|]�2ʐf������yh�52�r�!�&��*�B�y:��ec�h��=��W��� ��ߘ��u�l�yK�>ߓ�7�uA�G��i�%���C�����ڥRHڼ_X"�[s$�AcGĽq��<�t�k���2��|��H�UD���u�HS�z�5���9��^����=(X��e�y�!_F-ã���*��h�=`b����֚:җ=wYH���u��|��S�'�ʝ���
���<���h#��ۭ웧�j8ݳRj�}?��0�_���D	�L�a��X��Y�l Ҋӕy��/�|�B���Ph(g~".R��=M��d��=����R_����������p��.-���'����^?�I��A��_�ܕ�
KQ&p{ܘ9A`�i�7��Vᯠ���C�pwH�Xb��AY��!{T~��zU�CS[�m���X*y���s�<r��x��OU�	@�7�};x���'xɫ=+�h�I|Lw�;�y��e�J�$�+7�!vT/���$y�f����#��p�>g;�(�IF��Z��:w 3�uG#A2Є�<���2S�ܣ[�~W0C��`dp��l&�(8��t�w3�Ȳ�Te�����ZZ,iH���T�)T[�̪:��8�D% F%0���^	_�U�T)iNC�C_�fܿ�
�sk��ӵn�UAJ?�@7��U����l��By���`�n���-�a��ԣk���~N�u�����,տUiTe�X��F�xń���%�8�_E�̓�cQFԲ�;WEM^��m��r��g�W���:�%p`���1c�I�6�S H�}kUi��p�״_8���d@�}�"�^��fV���+�S��T���t6t@�0��`<o��������9A`����D,g	��=d��"2&c4�X1ndk�	0_J���Ze����lP���N���ҵ�w��9�r�����XxKr.0��cv������.p%����;���Z����XQd&SœX!����
�XG�/rs���2����Є�\(y�����Nߜw�