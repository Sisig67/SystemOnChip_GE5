��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���!<So���2��E�!�7���feI�R�34�F�\1uR�XO.P㤳��"����(W�����Y�us�'�V6g{���/�Y�^( ���Ne�[�����8�1��{SZ�k�eZɇ�FUHn�i!��Z�CZ���X�n��U�tr�Љ��������z]O������փ�=X�MG5�G����C��{����a�}�C�Z��b���>$�����z�[��l�;o ���'�����.���%�1k16oҦĘ>:���Ai2�L��������
n{Yt�n!������j�8`��Z>򴒈t�RJ�^FWwl�*�GR,�a[��>� q"��?SA�u��	P��A�t��A����}�R��Ѱ��ÿG�<�=fH��;��?(��ڞ���ăi6�-Yd�4�>���t��I�[օL؞�ܛ�ZN��<�����J�ds��#a�D؏f3�/ݕjEp3�ļ. (=�T�|� ��t��O���	Fo��8�05����a�{�,�-o]m�|q^�ᓉe�5H6��4�iU'��?��>�c��G�B���+���)�p�\��>�1��Yf�kn�0B��UR6�J.���{�I}*}��B6�X�tmi3 ��^�3�	��ݜ�T�e�h%�ʹ�&�#'�!E�!U9�<��o���q����W���T5�
%(�8���>#���~y��8�����t������iG�oI԰A�(���|6��vw�t�'����Z�р��IZq�Z�r�x&�|���L��A��Q��0���:��l�`���Z8<X^�I=~����F0
R��pȄ�֫p�|�I��B��6k���sI˱��)�6L�A�t��G �[l�8"6_%��NY�v	̚+Kh��7� ��%�+�(+������|�%r�������mO��Rշ;����>6��#��t����� �4)p]�3��� �Tʉ��5@��E�������ǃR�r��ё88���w�I$��h�NU w�'�*�G���h?�3�>΅�_�]�mr	�5��¯s�aA���w	��;��g��7��]kÚ��L�^���*�~�Y�艂�=宇�5�]Z��z苪')h(�9�OD���lUd��LͨFw��S/W�Y����z�,ES�?�ྩv�sj���Wy$��M�ѕ	Fs{���d�|zm�(ɲV��Ą���Ogu6���}�wV�V	��/vReεk%����� i:���0�b����^��s�\@�
tL��s#W�Ab��ު�xMyd�/8���lT��S&���O�=����$Z�+:r�*��9��|�ۭ���L�����\��K$u�1[��T5�,��m�_å-& 	�A�G42�^��O�L���,�����dO�b���$ �g�h��j����(_?9��G�r����Y,�Pr�%�X�i;F/jɦ��ϼB��'������'�3�k[��Y�+b �
�K)�%��i��۹RB�m�q|M���-�ZGA������gD�x������>�D��U��)#�K�G/W���JrD�$���c�[�d�֟��U�|b��-++���|V��EdPM��t�t{)��ʐG�r���ko�Tohu�RY�Y\���`V�p�:Y�E�fJ0/��J��Z�c7�����	R;��J!�����U���޲,��'R�n��8�(�Q��]bp{Q�d
�j�N�>׼�@h�Fh$�5W*OT�A59<b��U0l+���{�x���p��.�1=��}�f���F� rUד����	)/Ws��B:�!}9ۍ��>1,�W��ȫ)�J��϶}����K�x\}4w�d�L#�$�D��¼
B�
A������Q�tQ� ��,C�q�4�{��J�����8��G�CT)!�=�0����	 ���p��<H�x��}�x��8��qZ�q��������=F���;=�T�!u����PН���w��}����9��6�ґpP��@M�0�&B�)i�p���A���+&|�3Q J�X�˺��>�C�x�ˮnL_���o�D�??��5�'���|��rr "�����Iv�Ti`�l��=mbg^��\gE��z��f�}�=G����,Q j����"���tF��B�\�^ov(��u_��0����3RIT<�@:��!���{`�	�nu�,w0�� �_�%�SV��ѵzH}iFӴ+�o`�h���@19�>������8�}�X3D��ʒ��#��)P���<s\�\�tW��2�]<��Z����l��(2p;�kI����ikY��
�|�
DJ���(����KI��d��s�f������D ��2.Χ;�d1��e^�F(���!�'az����}SzT30�6!�,�U������7�s�-yK6��s���y�=1I��M��,�z#���8D�����+�g\��8��@�I�n�,V���
��1˱<j���˝f�[x��1�&"�`A�̒�#K���<ev:f)lG���pğ�|�׬Ȟ!��$8����泃�IͮCT�z;�/
ujQH�s�����U��+��[��?z���x���}���uzw�i�Y��[Tr.������)F�ZNa{�UIa�J�����>:��5��Nz���̟Ო�'���/�2�N1E�F����D
�\�����YjM�T�f�I�^��psEj�v�_��Il���f�4 ��H*�������."6ڲ	~\ڌ�զzu�x�m�
���Ϛ>�\��Ҧ/�ص�`�,L	�Ivx@v@|D�M��Z5�o����(���D�)�����| npV�)ƺjIB[@��5�����c&�u�PQZ�c��pȹZ7؃�Qr�X|��'=��#u��z4�P���.ߊ��c�_O��d=K��V���C�V�`�̦�g���: ׻�t�5����v����2p��;�!���,J�&S�n6���'�b�7i/�]�G�XŰQ�R��c�F�d�t��Tϸ9V�ͦ�K+g��1���n�҆qO9�&��9OG6����	�^.�;���.��!��$�j��6���p��x�VC��0\@����R"6�nuJ�<�~�`�j����R�(É����--�m}m�����,Ʌ����\��_:�^2"mۛv���F���d��흳��ِ�i��Sw4�\s���j=ԩ[�ڵr5����ʾ�TV�E��MeʣG��c�����;$!�����iY<G�G���� ̏��+�ȥ�!��v���5T8R�cX��O��w	d�0)|����Oi�P]�74K�d�qK��0�$Mq[�����2 ��4_�-�����|Ɍ����m�y,>]�[f�b )Eg?ز $Uh#�-���0V����̉�̼@+m�{�{œW��ps�F4(D�c�s:	���"%B��)��[�,�PZ�C������+�����T�]�y�>���#����$Ǹ��{f�-<���ˆ���s�6<U<Cv��J�U�Z��l�}( �R����UV�Q��
���<]����'�fhU���>�4."�/��;�v�p�8�~�PeɰWdYZ,�9�ki�\�r� X͗13[�\�7�$�M9șa_'�=vOa���Y�
���i�OqU�໺�����zJrq�m�1�'^���ސ�`*����GsD  ��H-�a	W켇�BQ�w�c����Q�]�3S�&� 	�P�p�\��s��(N�&�1G���*ML#��mn��j���'+N��W#���e'�z
wy�Je�sJo&v��C{įM�MT���)�`���-��KNs˖+��v< �D�S��ε�v��\�8&��ӯο�_�퓢�}�T��Nqo5�H�j��!lX|g�����K��������J���py��-�=~Nf(���W���\��a�C�k��̖`��h��[���*�	ű��1L˱Yɗv�"�V3�����2~-���3/27t)�:�
ݿWzXI���c���&��� un=�ϻb�g�UW�;|w��Kh5�A��Mb ;A�!��zď����������K+�O,)Z��\�."M�&!����!�Y"��F�P͍ �S�с-oom�A���#��H��m��?�0&���}$j#�x7�K��0�2�p�Z�Q�w���Z���b��!>i������bğ��p;	O)����
��Z�����7���w�W���願#~��D�<�@/�
x�y�h��21��MՃ�Qb�B�һFҸ��&8���������n����4u���yW5z�s�$O��~��t+:t q�eU���Uϣ4��u'`3��ꋶ�]����(�����y�GI�4�2+, ��|��`"���2�O	�x�[�B�-�LR+�,.pcs����������zc� I�$_8�טy&����+�K:ks�"#�5����ú�jr��>����n������lM�g&|����x���!X��'���N��S���<~H(m��m9Ȍ�nhMO7��2H'�2�pz1~�=y����͢b�0!�L�M�"Wl;Kd^t��nz�	3^39�,���忻�	��I��܌�6^i�V͂���$��.�U�I�����T>���)o���*��O7�#^s�TK|v�����\�~#~!�@��>�m8�� (�2�ɹV��������$>?����(7��,���a�c&�iXG�O�c��m���wtys{�6��枙�۬�i3*����w��n���gB�Ó��q~�CWuh�� �C���7-�i��3C�ww��@�
F��k��O��$������U���@9v��G�ym�wx�(���k3�+���|�G<�\]z<=pF3�FZ3s_~�~ahH�d/����z�D�i}l#�>ncHˬ�|���Z[�7H%C��_BG	M�v#@0�O�FY��#���s�r�U�F6��22�G+i,��rꨟ��y�e�|�Ω�wR�m��I�o�J�����Oj5��<Q.E:+p�L�Y�Ü�x���ū���g� ����.�G����XP����ێ�ԮD�8��""{p�a�\����٘#���Z�����5ҹ۪Ǘ�m�8��	�-$�$�!�X�2�dV8I�X>;�X4��߅��Y��PĠge�X�K=j�k�ƛO�G�AIp�����JHn5�n�Fu)E`�����T{k���H]�����K�xd���ὁ��j��7?~��,�f�m���>G�@��qm_�xaxG]	�9iY|�F��^�~���`�<D!����I�o���O�?l�:i�� ��W�'�Yc4���`4�r7Wxj�O�|��h���I����w��w����
=�,8a�]��aO��@��D��l��p=������k`fϘ=VHf���4�A?}���e��hH��;��Rw ���Żx��i8�մV8�U2v��`��^����ʕ�=-qj�p�ZW�X!b}�Q�}��*�C���/ `i�>�ь��Oj�V�����$'�����BV��g�9���}S�#}�3���N��.�Gy�WݎL�/{�l拪X���k�TZ>�J���-ސ���@W#�Ԅ����.����S|�7r�#��|��Y-R�z��Aw�A=Fz��Sf]wU:����{��mm�/�� Xr�Ge�v�^��H�L��a��Y��}��5����7P��q����X��T|oJ'mŰ6����%����L�I�/<�G( 8Ӕ��gk�9���J��d��I�'[�=���4����"�,�5�WB�}9��6aqU��:��4�ꗧ�&�r�s���O3B��;�e�;O�<ub]��L�X~afZ]�
9ed�T���a6��.�T�(��A�P���'��v����(��+̴0��AYN�3��@R�$E����y[6:����fj}�4��&}xuJ�ŏ���MH���R-�3�1�'�ꠧN���s�}e��178�Z0 �"�ٗ�`��	�������^&�
}=��w��j���.��@_��'�q���cЉ��X=��c¡�PJ��鵠�@��"�oEb�t>��UN{|nDo�3n��|��oʨ��o���	��	Em��t����4��+�̅�����HD9��\��?�?4��t�0���+5��x�1U��mS�?>��1\��~{Y��- a�:���%,���N�
UX��x�t�NZ:�w2���ƾ�Y�:U�x�&���A��˘��kP�u̅COt����o@�;�W6IFО>��- �P��������{�r]2��i�1g\oi3����'zBt�q�@��PY��|�X���T�Xw4�m �:��'��;^b�w�.�����G�XH@��¿����$���0�i�צK�g���7�A���#Gӗ1��GV���@� ̜�М����h�X������� tlJ�6�߆FeU���8t�p����R�����-e�+^�ڷ5�1�.R���hN�]�Gk
6��Kd��_��=
�0�P��KSu��B��m�а�Rgt������;��$$� �&9�ΎJD��;�~s��=2�KGoF�͙���"��?˝Ur�"�~}OE+*�F�6(�ل�YO�Â\1���YP�܌U��n�
�b��x��~c���d9�m$���!<�7��d����l:��A��a9c�-燤h�B�j��(�ț���LN��_��� �?KQ�B3�g�L�5FjD���̸ސq��h�����!"V��c������4T;P����y;]}��n>�R�=�:����D�3*;�lO�
��T~�rH7�4X<��"h�`sǲ�G�j;��>�����k��S��>��IK9
����,ZwC�`�b�*���5�Or�H�i8��c�����C��!��1TP���}^��LM@��u���y�m���zÎ@OɹG47�쓩�![0�������DO�N��
��҆<�ik����$��0��vC���ܯ9�a���*dl)Y��ϱR1Cq!H]��	���Ӥ�V��S�p�[���h���G�y�x7�Cy�\D&�5�l��Wk;Ji���Q��B`������H�Z�c��w�g���ڨ�jO���W���3�58՝Y~��h���X���,��d���9|��������F������3�);*)��p��u�E^��T�p.�h���S~8��<�?P�9a�Wݥ��԰Y}�t#�Lʐ�9R��Ο"̔P������]����tc=�����/U�3غu�E��A��A���p5�[��iK�Y�s�p�y3��h_���q�0��N���'�
��)��|�*J�^"%[��X5�?��Tcp�*���$�c�g��K;�~�'7)�+���sɿ7���uQ�2?�ʠ~X��8���t�^�l�����zN���و��$`R��R�29�W)�%���8����K�&m��pK�ܚ���u-�J�L1b1(BBB��%߾�����t�?�wZ�X�Y@�T�^�Po��[Dr�0��ē��h�#,�E����L!+vO|0d+��k��/Qܘ�y���sǵ�`T�Map����H��Wu`ˆ�k�,�q4ߥ�	�Ц��P�*���Ǟ���<H�ZJ�����i�ЂI�e T��		���*y�fH:�C����p�(�>���0��6W�ŭ��5�y5gxPHa$�;T�,D�OHH�'Ҁ�g��]�8�1eŧյ��чR�/�.������Z���,&���E#��&��l0��T����w@��d?R��|�>���*�s�6�J��@J/�ߖ���;��p����C
x�$��iX����i�qp��ʇUs��&ӵE ����DE�<�����N&?��G�s{G2����[�@$�1�̓�3��e�;�FoC��K�D�����<������U�j�]�̰�- h���^�Lu��;�}�@%�thA'�-I��h��=��*��e���]�
�3�P�LW��`��DS���rx*��5��(����P]�/>����c��F��~�d��RxƁ3���<����ۣɕ��GL�E���~!������^Y5H7"�����l��g��*w)��EN+�E��fN}t��pi�+�
�#0/e-��5=���r,3L��?���%�`����aʑ�mx�P�IoLN��8̙�?a��*�� [����Fa��pDj���o3�\q����5�C�Go|�[ߠ��v��<��� e�ƙ ��&�0�qZ.��R��Or+� �Ue��1%\b-����J�����q +;n�/p�ݠ��v�Db�o�i��ϔ�|��^�!��Dw���#�L�l�<y%_���s�t� �����l����╫B����1-ޟ���ӛ(Q�m��Ѝ��#Z�Yg�E���,/ ��"��	Ïw~��oynQ4H��[�����_�ř� =vv��W9���>&�.I�Cʛ�{e{KH�>�S7Y*�� �)��i�N~Η�# �O��Nw���lU�)ۦ]{ڛH�,= �Sسa�rz��4R��1�>7Xps5Z9?V'Z�(���-��w}/t�ܻn�u�����zO��'X<TM	�a��|۴p����^'�L����2����H�ac-F��X�q���u㔔
����R#_!*���a~��m�f(����M	y��m4�&�oK�w����J���By@qZ��1S�>����6�.R&s��u����2�[��Q�\9��c�F��-dUlsez�<��"�ʳ�l_0*�VʗԃM��H�Y�Zg�����ɩ BF4r���H���I����T�1��ܿ�.V���h�0�цA>�����7�jN��X�J�*fJw�m�����ʑ=]���(�\B�j�p��L~꒟"���t�=W�aVr�"CR�5ˋ�����z������J������U�!��O��>�O�P-��$] �_-\{,��R�>�S����Ybx�*]�/�<�71&u����%:(��cC�uN�d�����ҖK�5�q4٩����J���<�_><c�CFC��v���W�E�2������ōsE�jVHO�?��<�mC�: >@��U&Ȭ�֭Ë́X��;.�I�0!�j�)R�p���+�Ǔ=bۄ?��������UY/�0-��L�)�>l����zQ���S=�~�ֆ���a�ʦ��]��y�X6�\̐xIwC���8���т2�)����4���v.A��f�H�tyGB1�u��;.K��\P�P���ɓC6 '͑O���� .?�����4��8�>�'�?�n�^��K	��9�����^���ȝЦ���K?��BSn�mt����<�"W
1�JIWK�.��v���<�ɯ��*x��Qv|%!���(A�~�ԭ ��!��&�#\���!�� �������4�$fJ���˨uԃ8�=��y�ѾY=-��|7H�0�9�,wJq��(E����s�~��V�
`B���=�! %|6���l�����soT߹�~.	w=��th�	������HU������}z���g�.dZ�t��2%��5�ɭ�E3	w�t�����}���e��`�����Bk���s�X�v⨾l�:�(�Q�_졂�{��کK�YoJ�d�7-�q-�A�굲��.�	�#!_��["�ES[B�U�'���쾬`Vׄߦv��ϓ�,�ĤO!`�`LP��uC�s��%�%�Q��/�׻������8���|���PI��j��|��)�M	: ����2e�\�x�fi�o�����{Ht��������[:�x��d�࿰G����Du��[9'� T1�1<27����R.��FL)����
�*Ǿ�=��\�7H*8�5�b� �K���$U����n��Ro�~�y���V�XTbD,����~2#��P�%�wd�w5R�
�<h�(��y��y��gr�l?�FZ��Ej��6���U}�����
��Ŝ:_�kx*�e,�p=�[v���$�@�$���k�US���t]�r'�
�YH���|��B�)����-���i��0<AUe���`MFE���ݎ����]U��n|馽X�7Ii0Hu�괢#��M8q�; �@'����1C" �>���{���&�u֗KH#J2N�t�����9�pD�S����b[�"���.�,�ptנ��5�A�g�q�Oמ��c�
�<��������~ܕ����ɻ�65�2�� i�Z��Ed���ť���ۙ�&>�]�t���ܝ4�s�>֢b����oQ3�t��~]����0��-
a>��]�dl��,���M��������@������=��j�&|�u�)�O���X�nr����X^t}���k�dE���
��S�{��h���ir~t@�iNt	�*���5���?;����%����j��gu6k��В}W��	�tܢ��uW�f*r;f�	eoq��y}m
�h����ƍ�RM䰏�_=]\�U���q�T0�:pS^WF��򠐄�gf�Ϝ�H�?O̚�J��RvsҥG������J��b��b/;=�٫�57�Xn��}T~l���Mѥ<{��oSؙ���i�@qb˸�=�("i�9ל�����}�k�j�d��/X��z� 4S�ة�\�Z��~��MI}���c�`)w���eK�,��}������K��5Z��N
�px�v��T�RƬ�&�`s�L];����
�u���%�[z�*�gz�6�4�@o�N������;;��!���ۆ��dx�N�Mh�dj�a����ڞn�&���J���NPy��B��1��Ú��)�
 �?��!�"Z�������~�XQc��r`�]X=X�j���O"���#O6����oE�8�&��i�:lޤ��=N6d4�M]��\9KsC�>�jG-����?c�7"<�e1�R�Y�dF=�c�Jiy?��~�sk��6���c�����2@���*��خkl���f� ���YInӱ�t�$�u@�h�!�v� y@X�Է�ح�D!Sܶ3T��l%&1V-I�5�͎�P�58R�c^|��_����W�^(��ʪX�;�i��3�u�����QK�����. m�=��ˍ��Q��{I����[��@��b�\�ae�}��;�W��N���Ht2���9��qAX� ��˔5�T�bԋӔ�7}�=�O_,��at2�&�<`�ࡈ!��;��\�Y�#-����}'�{�Pta�D�$w��I?�=�'ľ���1�<�L��3R�; (�Z��'>J	�q�ޜ^Z7/l��$R�B9k�W��׌��;�s������i�[@ ��a�cٜ���|�,17��0>G+-����c:DT:�.t�,Gl6���>�S!��W�r®�B���_��0t��WI���`2��ϡ����V+<���Ԃi�<+���kҀW>"D�X݃t�A��<�aʅ�)�������ǩ�wM*ʦE!U�{_͓btp���"�)2�yu�V�2�EHJ]�'RD$(��6�=Ea�ז��K���j.9�6�P������Oʷ��dUv�/�p�a�l�J�}����X��@�ם��4d�z���d}�����u��U���K�D'�[��i���\�vO�|���ñ���6���6J	��O��#9�8R-\ZwR�r{hpUT�K�pk���\G�]nf
'�j4�9�:��1ޫ��K�&Uh%�׵e��D�I�F�U�e�ĭu�g:���\�R�^���"��D��]�p|_�>�M��.�&�ˇ)��L�όa����Z_,��AY�s=&��n�
�ech�(�U��.a�$��1���LZ��H�@5�=	q1����L�^�y9ݴ�U�<qC��I�8�*v�����=�J��7���e(�0��
V�?���P����J�4�C(ua��]nk2H�/u��r���L��������U�D.k�22E��[^&F.�W(![{�f2���� a%U�F�^���K��[�>�@�.�5
�ۍS���(��M��(K�L�+�;��}3�ڍ%n��7�T�v:h�ᙴ��{ld�z6����S���&���ƹ�����\���Nz��|:�֏���T�tw��!�@�FHE���R@FX9)��N�rP4���Q�ep8��7���y��ۊ)D$�-K�W��bX&t3��.��8�m��9��w���-��={TQ�H9�[��]�'rfȑ�¬ҩ7�U�Q��Sog:\4u1�Ķ�ܬ�����l���E��Ӗ�S�&_U�s�������������q�Aq�����~~й�X�K��_{�z<���L{ �n�1~��E����$/�٧�@���Q��`��[ ���b��%X��bw[#W9ڗB��>�A�Li��i��s�\��pg1J!bk�?MT�=,� �.x
\v��uA[%o>nY��x�-~�1�����5�4�*��&K��7��	��E�_���6��a~׾ca/�0R{�;��j�W�K��W� w�,�^r$�{�n��A٣wDP(�i�t�z�4�}HR�ru�}ݖy�Z_t�MU,U���-E�GK��V(z����]-ȴ���mg��{1��",ߙ�e��tp���/vy�O��놺+�ё��`_�E�mL!��*�+RW_^נ��w��b3zy� ~�ǟz2_^l���ܤJ�7j��
U�ss[��Le��mk�ZwVYR����&B\���㒊&lUc��A%�Q��\#�V�vj�%�Up�Fә��iRk~��i�%����>��Ϙߝ�.�'���V���xsd'�ҫ[#̾�~��p/,���?��"~�B*cz�6cm�n�a a�XI�}�~�����֐C�'��+�<&�#`�s	�7!�K�Ҩ�	Z�x�S�lU�W��5�T(XM�R�]�y!���������]R���rdu3���Gk��o�D�M�W1x���y��Ů��lmC\�?���nc�ӻ{a���	p�	�[��!��<�vz�&1Ԑͥ �9T�b�|�6�����LUtڌ�>;��R=�@f�dŃ�v�X�!�fh6���<;inBY��=n���e���R��4����l�S�9���;��qdn:^q� /�_��r\$gK���yYDS<?m�0�F�$o�W	*LXIVb;�8GR���SR�v�T7r�ҧ:!����^G�a��$۸��@9���`e��^�m+��/�JU��&)�B��̵Y���o(A����!ِ+�4?]{}�i��.��� ��,��Yj2�l?�������: �\7����wa�j]ɐ�"~�U��&\�W��m���5ol
�O��i�����*h����m9��}��Hv���T:_[�Kk�
�hg�_Q��:��+=#�]]p� ���k|=�粆A�x����F���|{��l�M���
`,ʸ.��}%p������	o�p�0�"�hAG��u�ل��o�L9�ϴ7�:}M)/ Z����d8���$�
r��B)�#uU��ܰ�Y�p�Ka�P�3ޛ�fB��E5��H��e�(�Ҵ�U�	�ἇ2�x#�Gϫ`�됱D�Z�TU���������:S�׋�uO)7a�U�Ͳ��)�٬B����Ɂe^�Б�1.|�DA���IL��4�Y=܏1�5��3x�J	X<��GH����h���22���jB��ֿ��䒽D�a�h�I�E?]��և)RbNc11�)�<G�ޫ�L���N��ʿ���6*����ӏ���&\���h���������,2��v4bȩ�����*QR��}x�R#K{�GV�?�����.h��6 Ԃ�JI!�;���M��V���ue^�O��Dl�BY	o�o�Qc�e�Ż��$�"�$��j�����(��B{dc������B�9���iH�o�d�z �xIi���k������J�ZA����J�H�yǽ0�D�B`��M>yߔ�L�,)�ۈ8i�V��Q��<{S%Hy� �Ck��%��N��^N_��Z�Qcd�B2�K�NW&�ޭ�
��,������s��sb��x����~�G�ρ�n'��K-�_�e>JY���c�?m������D��HI1�I�O=BP�v�آ1��ύ;��jҢ�`��W�3������w��ϡ�s���3.Z�4��-tc0@�Q>�޻��L�ý�H�F�,���w1-���Y&�<�r���WQ�L�I��w���ַ�	v�r.X^���tj��s�	��B�\�����d:2=|Uq�u�_)`lG�",|��؛��e���Mw��"��.ê<U9.���%-ȪK 8|�8L�1�}�`�$�g����b�����.l��V�7䠣���  f�����T��{���P�kQ r��j�E���QkS�jC,�P�W���-�/M=]~�g�a�|�|a�F���7�hy�h�R�PYCN�4�C֋�z�N$n^��M�H��"$�Nz�>ϋ�c�3��fv�u�2��\�!��LLn�@]H�COg_-vd�:�N��Ҳ��CN�7�ߺh�zZ�#:�x� ����G�6���[�s�1k!E�!�.y�F��<�9@�0�O��TJ�d�}*�1&�==q^�w�X�+�ja�����+���D���}��|$�Yqp;�쒁��ȵ	vݣ�Ea����6d��2���}�_�(�͞b<R�D���HjZ��ѰF/uK����[�G�Ƀ;Kծvg�BDEv�=���X�>��'�����-eR��!��cѓF����4*�o��I�}���[��/F��n�N�`�����b��5�.��i0�����PyYZ�h:���*�z��q�y6K����<;��4�}72oPא��\���:�V�PT)�AwJ�U��"
q�>�0�]�g��1�.�じ���c��J,�~	W
�-m.2
�Qwo�b'�1���-�(>�੓�m��$m>���5;�澾��5mn�g1 ^X��DO�W�%�	+�O��nC����-�Βͫ'T���W�:��'SP=�z���pp��7��z��!���,����]^ѷ��&~SB�F��R9�|����_G��WG%,5:���� Z��a�&:�5W�Y����=�Gz�tr;��1b���ӷK�ϣւ��>̳	9��[��;P֨�/4`Ax6�ؘ�s��\]�Ny�)w�@]|�`��x[��uI�]&�[��6F=3�~n�wn�ZI�ώ�h�q?�Ⱦt�"�5���d�(sܖꘐ4�� �*X^&$��.R���$|AM;$]�Jl ӊY�φ�e���D^y�V����x6|0LB�3�k�`+σ13Q`�c8-'�a�g�jp�����:�����?�	=���7�ň���eo���n���ơ&e���M"Q��*t�AƐ�ݱ&	 ��a2��v��w��>|@�#}�M43$�h�6Ӌ祃��ޢ��K~�zŎׄ���@d��b����w���4� ��Aգ,Z�}��{b�D���#Q�YV׿�/�A��d��jP��])�h=����~����G�} Qa���o3A� �ҪG�;��������[f�s]l��$��hƼ˶PǦC��i�O�y�y����_y���#0g[*���d��G��KI�.�����I��8e�u�[�m�V%!ȵ��O�zz�w��ܧ��ݫ�y����=��)2ty�q�D��͒�C���zX�^"M�u���|,8�w.��Rk���K8��?a������F(5_nU���63FQ����<ܵ�aX�Ym��O��q�Ս��P�:I�������i�	1$�	^_vp ���,���5��;O>���<�^����OխAM S<���?��%�b�6��9��s�}T:q��.��N��eD�/��+��	G4$������$�����e~��B�h��YD�r��q���h��Y�2��ك
&���p�}���u6�_���<"�|h�,�?�p�e�U�p�ˢ��2`.�"{�Q|�ib7Pp���Ak�C�$�Ơ�밪���@������䎥s
�8a�a{�ܼ�Ǟ:�
 �������.�[𥕃c�T�����%�J	��r�wF��8�A��;g5\���ǁ,O�&$_�bƁ�TK�>*�u��q�%�8�o	��he�~e-V\~g�M�3�j����S�G �o��8�F��;���0L`-�Yؗ<fC/\8Y_��w�U+k.g�L5|2�P�����S
�~T���'I��*��2I3"�{vsQ~ Y�������UIvv{��~�8Z]o|���WЯ	��+�x?�D���5xi�X��1�h�|ZM_g,!�vĆ+���quN�����~Jw�e�\��������-J�޷+�dH�nh��d��HI��+��Q������o�D�rOx�X9}�f��ש�é�%e����zL���Me�N%ƥ��d��$�UY���U�\����:%�
ϥ�e�!�ϱ�9��HiYp�����6^7h�[�s��fkԟ��¸�)�:����C	S�}���Cc�?&�a�G�m��>���1�B�S^� �p��` ��g��i�b`8������~�++}�	~6���X&u,���zNۭ6j�n�Nn?m�P�)e"�*"A�(�����.T!4��N�9�$���Y�	�,I�	�y57$�x/������K����l�
k��LYM�>snUˡr����$G���z��.1l"�Lo�7������]��rFg�4�����7?���i��mZ���@lN�Kǎ'��'��BI�yy�!�7����z���v�iv��� ��N��x-r3>Us���e��4����w�i�\��9Jn�%�B�B���a�9�/�?��~G�֑�9�l���;e�;�A�A�R��ݤK�#׸BM���;�K�!�]M\���PH����X���f�`��r�����|�\��F?�Il��8|>������D��y.��!X��Y��(�em�Ve��1����6B\!y��t�Óđ	�� ���'N�t�u[m�V}���;���D��tE�O��F���zX�jꊉS ��� ���R�$:�Q��L�(�f S��e|GO0n�hS1��W��3z;��#�ꦛ:������K����[ۛb09��#�E�1�G��~�kK:� ד���@\!��a���5��ə�:��nO�mb.��WU�Ф��;���h���JU'=�l�o��=YC^t��֯��/� �?!���P�VٰV:� Ŧ��2�3�FW��Y�魯�c�# d��n%�����pխ�r�:X(5����ix*��z6�E���z.�l�\%���7����{TN7
)�f�n�� &$u�,�P��O<�G��)(�Z������{�g����[ �
�+��@���t���_:m۾K�0�oӀ����կ��z��L�1^~G�0��^72[����{���Ԩ��m��+�Cr���f���_A��少UX򥝹��Ū�8*�i<@�Z��uU�j_H&�w9��u��>��[���\ʧ�y���4�ZF�&��3�ۿD_|����^���)\�c9�F��z����*����x��':�+������!^�~�.r��C0��MU��42p!�p�u�&^��Q>�9L�Cn?���Fs3^���={~��Jg�I�R�[���N��e����[�9�##��Y������`�\��[F�� e�:����z�H��1�(rAA׷b�� @^
7�s;�ۛԥH_�JhF�ca!anr2
6��w�Mw!z���25͒�-qޜ���쾃DZ�e�t4���� �/D��8�ˁ�߈N�$P�D'�P�I�	y��L�f,rp#O�T��r^����2Lo��$�#����I��sY-�-�.�=D��cl��ٵ*ν/jhnX��N�*4����F�L���#�h0�Ľ�	�p�����Gmfȷ$�áf�V������[f�ʏ��Ӱ����>����v G�[!�B�t: �C�.� � �'�U]��[�iO^�K���w��n������>s�q�ꈧ�|
��b2]wl��p~�;��\�,�A!�3�O�:b�sd1��Bxb�͐�j�	�v�[�^y�7�W{�,'K���۟����[������p`<U�;$K@FQH�?��͠G���'�O����)hh�8d�J��_��7��0�sq,�ߎ'8�8G���r>Z3n�. ko`#�oL��OK�+��R�ñ�4�8 ݮ�M��S4��P5��ķ�� 'P����(�V`kUlS��Y��oxS>��V�Ӱ�,p[�n�"�H]�/
�����W#v،Y'~{�����$2�;�����R�-�u���
+bpt[Ǧ+�Q9%6�V�q��KCV�탌�_O�t���;+�Y_����&�uý"�&�ҩɩYY�i���.SB���MX��[��hZ��F��R��X��(Ξel�l�9��{�|ee*.��{l(E�KEj�f$�����ŵ3[�6+e��l�V'�9����M��,yv!C$<���Tx>ő
|�VD)���H�;��	I�ӈ�����Qd,�_���vlT_�Q�$�=��<��^���G-AZ�Ib�����p�+ g=��<��Ă{AD��%��t�H|�\Uʖ�q���V�@u�bM���wV�A���
�� �;�>�"��̲���J!)5/
-h�����9�F�]3�s�����zs߸��{��
k��aE�ނ��׫����WM ���j�gkR\(u�(�;�;��X|�F�����C����0$���m���+R$/�'�91�P 9��.V��۲�K>�]H�ԽT {2�Y������&�z+��,��v6� X�K8��,�o�/v���OHn&N�>�_���ݷ)m!'C�z�R$���zFܸIȏ�'�o4�hwBsT/>��}����@Qꨎ�Rꃹ�h�e9"]�Z�$�N�bM��7HL!=M=^<���y9BR�Q͒+,�4�������ԙ�o�����)��������A�͝��$-��O���_�|�tα�@q&iV:8����z���c<�LN9�e2�Ôno��������=�.��@�<�W������)Q�=蘓yq5wE�"I���`s[�*�5w���ɐ�k.CHk�_EZ��/�W#�y1O��leWՋ2L�66��>�J�֧Ħ�-�*�h(DTE�n�V��N{�4��G�����[V�l��N��~l7�/,��9���o�����B�#�l�����v��^��O����Dph��:u���#L����X��x��YPxt�|�;�ģ�0o��.�RD�̸a�l?�ag�ll�%Q˔��eocV�)C����|鎓�{1OV2� ��cW%S��[�V�p�Nn���>�#,�ͽ:w���a{�0� �R�E�?������<�x)'ӱ>�P�T�G"x�#���&
�JF3C�Z�0^�pALC���nn��,hזN� �����}C-�Q~�/R2�豩�kaGi��ѐ.ˉ��w��N�ɉ���Yĩ�FȎs@�ӄ'	D ��
�O�%C*ͽU;�x�mB�X�"�D�8�	���g�ABԨ����qw�e�`ȯ#�sd��Y�L���yQcX�2#�&2�\|�-�&�%8ٰ�Г�)2o%+s��chC�YE�Js�~�G_%�p�')�&�^��P��o�	��@�|l���y}��&.z��M������V�	m�����ynK��"#�[�}f�P�����ss�{���4�f2�6�J�����jx���ܟ{���[��nn�6����sr-�/�I-���z��7�*A_��soH�;�}\~K$#B��}�8�B��u8*y4ʣ����B{���Ov�YrF:��'���p$O<%59�GA��۴�L�����t�����?u���)�Ƥ����*�T�ȼ���s�N %5ɍ���1���a<�z<��|	�9��[,�D��#t#i���{=̴�8��~��E�هS��	�A��Jz��Y8���p�%� KA�a��@�����<�?�A�������b�N"��11��*w��j��/��Ã��)8�s��������t�^o��O2��Ѩ�+�bUg]O��U�V&�~��|8�+߈�5#q<�)�&��Q�Y)�/��!�_#*���#��r�<�\�V��[H��t��;$i����9�`mKT첲��b()b��R,��޹syj�~{�/D�x]�b�90r�xڕ�cl)��GI
�^Y�99����)Bvs�fHٲꃨ�N�ȿ��W�C�#��6���C��+�EB�$!Q��W^1�q�������X]Қ���،���Q�"�}�ru�gi��l��drWU-w�Y�=�zҽ��b��S ����}g��z
� �a��0Y�;<�Oԫ�=Z[s0��C��&�4��daۃ(��2w��b4\��|foΜ=�?;4 �y@�P�䝇t�ܣ{����Z!��#m�_	%�w���$��σ�%�b��1 ?��r��v��y�HSY���L;\5Ok���ZrZ|�X��T�H�W�J
��F
�$H�уN��:��&�n烮����T�e*��{�:��`�оI��.bK�c��S	� ]���Թ�$2ƚ(jՂxS�|[��)Q�2
x�7�e��Q�wT� ��� }���9�"�ԇ:a�o'	a��sԓ��SI�-����j���}��[_h�߫�.}��- ���������+fmś�R*A�ݩ��17{�Fo�(u�H����M�_|ƕk�IP���K?b� ��������,�V ��l#��<�Rz4	�����Q!IΠ������
a�[�G�U��U�ɖ�q��Ƀc�m��&���+��+]?��K#*��#�,��]��Ia8�
z���syB�j���y��eG-��x��_� '�7��q��*g��?A\0�3ݸ����	��H�Q��k�wv�s�a�x7�ogo-j��r	W��F%��I�\��V�
��T�M����3q�� ߴ���c��CEZA�� �wxI�����NC�c褊̃���"���$��
�>��$E3���^�����CC��s�/@��W/?Ȃ{<�����]:b��3��K5A�QU �������e�	7�ْ��0hd��1U�W�H��"��	�+�|��wi��[��TA��!?�q`��ܽ��o~��Ӆ^�I�V�*L>`�C�z�1��T�c2�Z�H$�o��2�u�ab�\�`�� X׾�&�ux5B<9j�<�� �`�(�c=�����J&8�\hU���J<?;��f�
X��nz�D�p�b36
�`�V[��b���qţT �C"@�i��S��3��k�'�sӀ��Ug7N��.�|c��Y��^c�f{��-�]��Ԣ�ڔ(��r,��nY�ߴn־��^
��{�"����FC�C!�vt�o%��I'������n�BaQ��b��rP�~��D�u�*��y��0��I��X)]�\����Pf���N�e�<]�}�Q0a�j8��#�`�N�w��L������[�a&���!�� �C7!	�ֳ$7�w��͐>gZ�U�Qf.a*%�l��;�_�|�b08 ����tUlR<!BU�l��z���}yU��"J�׻i��Z�3jo���>~Z�<����c�O 6"OͦI�ي�\��s��`}���r%�Rݫ�v�
����j���Sw��B(�sdԃ9ءQ���W���Z��Ja����f�Z��H��4W��JB�Vo2&.�i�z�Uo`�K���T��bua�b��g~+�k�L�)o[�k��^f��m;��r�<�~��<|�t2F���a�?�O�}�a�A�@>�bkU]��P����@�����ڛ�ܳ b�M���KR'y���S�;2��=��5��h�b5`�3�qW���R�n4����yQE:�I�>0�ީ|"ĪЃ�������uE�v�fU�$��2��5h�:uR���,B�����h4��E�RL��T~D�*X�!cp����a�etnD�1��U���4��L�&�� v�0����mV��*���� ���g8�<��R�ʝ�(x�͞ݛs�C XӴA�����L�	��޾�7��>�<��j���lE��.;c� ��$2-�Hf�E;��8����g�!��}2������Lsy1�ͱ �,P�	�����Ѥ�����ip<ق�ۿ��qׇ����/�8�7�OC�N��:�ɿ+���«L�B��?���?����w��B�o���8��Z�*H*d�u���i���!����"��R�j��l�v� x����dA1���T�mk�M�t��m�ߎ��/�}�S���?m����BR"���|��t��w���MW�ec��
�nwv`��$�8��K(i�X��+f�cǃ�f�w(�>@|�1>���B��[5�Sj{���*�#�W��햶7�Yu���Ʉz�⭳�ٺ�-)V��=u���0����]����氁<�Fܼ]	�k<r��#4��M�� �'�8r���_	�ܷ��gy��*�J�ĉ���X�%͌j��� �W��D�N6��W���4�;>�u�g^w�q?�M��`v���Dph:Ù��V�Q�)ܥ�����T�=��MC���gu	�����a���n�`N+���7�K�1N2�Ȏ�~�
Y_�k�qV�:��d��E)e��@/0i�m�H�_VLc���G 	�=4��?�kG��	�#1s>7i���q{��m��������?}������7!M�a>7Vvqe(*��T;Y�ۍ1AQt(!��얋�_Q�ݽ���A��\B���ئPy��{�O>��
{[f�L����j���6��X6!�����8�8ٜ�X�[��ƒ�r֡�'��@9�x 	�k��o�D��{͹���􊳺��r_���QVX��T�$�[ w�@>P����j�HGZ�(쭔����3�e��Ύ��4Ϲp�}��?��<w
�O-���b�۰/\̼IH�i������t$�J+.�gg�x��@l~��CRĭ��oJ��㢍w⦁�Pk1�7h582	�s����[?y��Tm�o�l�d!�M/��lXB�N���N����QG���j�FM��3�eLR:�6ćuD���s��7b���xj�"��?ޗ�&��MQ�~jlv�G�%�d��= m�?O�a�(~��2M6"T-�gs�'B����}��4�K5�_�:=�D� o(V%��d��N)7{���q��{�Ե���� 9���1O��k^&�ȣ��Sӈ���,j�#�cB�v~���"Ǿ�_*X]���ލ������>tI\F��iϛ�)簻�~�o�z2͐�g�_˞����1��j�U_��n�#��. >r��"��HႫ�Im�0 0s�ғǦ����ň�Uӳ6�������m���gN���0#�-����P@��,���<0�����.�FF�V\d�~(��s��@�h\ܲ6�v�y�z#�N���b'�~%ɂ���'Q�/̰N�/'ԅ��b����S���?�4�/��@����0�{=,���0x͞Y�>��O��u����PA>�8��A����"ĳ�������|�ς�z�_`p�d�)ì��AcIk�'zL\�F�>P���a*�$W2��?1��4n�`;�Y��|�LM�E �֣�	�_�_
V�	�Z�#��:&��jBy��u�ő<�P�pA�4��Ojvn)}}�n�4B�^3#a7lѢ_�,��j	���û�4�<���, ,�A��Dxt��S���_�f�$;	Ŋ�#����]3���O�
A�U����[����+�F%a��<m-��r_��`n7(_� ��j���z�B��a�Du�;
��-�]������}�,��%��|Ç/W����g\|}�S���$z��V��n��Ʃ �wA+x�":#���Y)*5��\w�F�d�L��J�����/�[�Z�׃��A���G�����m�7��Y���-����R�!xH�WO�ˢpg�=b2�e�mV��it���Ûkļo�װ�����W��f����#Y���]l��UP;�owT*瀧�Ya�D���fr�38�<��9S.��`�]*�c�Ͳ�qVJ7ΤF� ��J�:^*����˜HT�?�����I���o$ ?X��GL�,��q�^OQ�^=�����c6p�^���
�r�'���W4����:�;S���@žgR�5��%#AU�"��>��	w`��M��&��G��LJ�u��37e�T�I_�.�v�D��>jE������%���8���������ig��Ē ��W#�x�9�z2	�\ ����m�m�v�[CnuP�i�9���K8+�����`�ힿv��Oն"h��?*D��+A�Je���rP����d�����:Ԧ����h��d����eQ��'�e� �.�Vb���b>2�-��bZ���%���<B��g;Grr�lE�F��d�/!L\��^jM�PH�|{�	�+�:��c~J,V/0��n<���OӖ���?]���k>c`���	��qUb_��sja/(�2�NOD�7��[��,�>���ץ`KW0������f�ɍ'�׾����ە�֬�r�'Mp��n�yٖ^���A����.�����"!O��jϵ��A9xNldU�{&˓��+~�xt��4�LA/�~��iA��2�U���޳x ���ӓ�AT���C.?�oj��K�]{Lml�O ��O�d
�0��hb�S$�-�+k�U+�h�ECRp�|��}.E�j������n�H�dpp��s?���&�w��˦{2>;��������7`0~|7͈�
@��,�g*:\��<�0b�Te�T�dX�* Cf�� ��B�`���s��"Z�x���N�0d�6ܵXL^4P��N�	�s���^�{����K򦬴%�D-ӝ̥���;U{������#�!X�s�@�1G��xܬ)���(�~�p�SH���;UWR����^�@&�D9a毌��>ƂF�����D7�������͠���J�(ؒ�_A0�7*ê���	JDe��b�5|Y|�@`w�3ꙆB�|��D\Y�~�w|�]nq�y�m#��l�X���`��a=��G6�"7.e?|�x��6�iM�X�L���=�hy�;Bo��^a���#��Y�wRP6xҎ�1�ln��K�t��7b��v�T7ڿt2�و�7g�z�8�f͟r,���S�Ŧ�lf���9����fh�ݼ��~��ʓoߐBf�*t s�c��:M8��Ϸ�2��N^�`���^D�� ,!��88,v�0��m���� |obHq-=c]�ɑn�hb5���nx�٫k;��4��UJ�O/�5�k;�	�:@�P\{0\��aY�d>r�3�������=|�U�B7n>W�f�߸���s��e���H���s��ԥ��5���i��M{8��U��ܙn�����)�)�_����^k���Gf��S�p�Q\BM�d�r���T���ȧ���ѫ�i�!閭��Z�6h�m"
�|�!��/H=�\�w�Bm}��&�ju*��\���L���o8���o�B�=K��3�_��쬸�0l\��^0:�/���^���a�����{H�V& ��y���uYi5���vV�d��rv���o�M�((W��?w�i�q�����H���֡��
�<W���V�k����C�?r�;Ҝ�<��Q�lG�A��uD|��R�d�!Fs$�3	Dl)�FP'�׍ӷK��Žt�Ҧ�Q"�+pU�ąm�;�V�3d�D�􂇎�țj��D#����,B�����֠<5��|�\��c�����P.4/��Dކ�����L��|L�vϕ"@��$ �N��0�+M�k�9�)x��!�h`V8+.Q�����h�e��0���A/o��$��j�ft	�x-nj���HŲ�����byj@��	���\����1�;D�)�b�{�>�!#|L��2�s�_���<]8��t��p�tk8*`.o=⚧�{?VZ(</Q�a���닮zg��SVۺ���I�|��#J��)�<;\���T�\�8��pQ��x�Eoͳ
c�lª�(΁�(0 ��_��D�	NJ0�$rZ��O�,�Pbw86�����Q�-5!�rI�n&UsM�sd��̖.��/w���;z�[$thjkڸ������5�p(-�}�C��KF�^M�G���[f�Kx�gN��da_v״��l�L�v���}Kv^B��H׳�n&��J(��,�D�堮}��F
�v]������Ɂa�+�fXY=�����դg�W#_q�A2�6o��B������c�� R�)�1�b_��#����S�g �@�Ҁ�5�̈��沖���`|!V>�M?\� ���o }B�z���5���8����!kĥP���I�Nf�m�et����;<��.��Ш��8,��Ѵ�X\R�?�}E[:=��HY�_9ΒdEj��)�_�O
ȴ�k�/�k�ԖF� M'�5>��ME�n����� p{)�����DYܰ��v�b�_t�g����ў������w����Z<ǋN2 "#���f����C�4�m}����ulBigx1��@���[���YW�0(m��-i].�T#�rx@,�Ωs	"sܠ`�L!+�=�V��[!��~ݽ=\;YD��˔Xt@?mMS�D�'��UV���2{Oۄ[�UM>��i�v�m{�)�!d�� .���?��&�.�MտE�@H�({ܩ2�NM�hߡ��qD�sj�-���LEqc��\�nT0R&,�rjd����$\�;���갟;���g�6ܮC�,*�]C��)��3��yJTّ*0~:'�����rSi<�p�vEXd��C0lU2 'ǜ��(��x .�ݭ�P��c�f��ްd| t[�~��<2�<@62.lZ�)�>��]�Bu�j��;�Tk�IZ������N���62 ;H��{*��4N�3��Z4x%Xh1��^�a)C�	8��5!B�'��Q��������+����-D�Uۘ�ίK~���p(�B^ƨ�r;+��T��q5���@?^ǽ�)�'�����p���̅�1J�����#���n�������N	�$i�ͭ�~{'4db:]�X4�� L�S<;�%��C�a9�+�g;�����9�j�d�q�S��N�$UI�e!=p�?��y�}+<��EE�s�Xlz���e71��l������M���n���:a8ʂi� �/���[��ؼ�@ �)�h���4֧��3��dwCX{z�Y"j�մ�@{P)���.�v�?���`ݻA�{YT�P��d����'SJ ���|Q.��J�|�F�9��#߯?<�Y�K-�
Ɠ����rE���üٞ�/�R	��.�z%�yЩ[��Tu�-���w�(NX��E9�FOtA�3���}}x[�D��g3���Vww�,C�/�Q��f�8����3JAr�{�A�<��&.���G��駫T�L�������9����cx��q�Jx���bb"<it?�|���g��>�^�1����V
���ͷ�*������a��8bݒ��6��֡x��\��(�CQ.l��W��� SVK��gA̐� ��|	�{E��nw"ۋ�>l�T�tg?j{�o�a�?���1n@��,k���H���P�Q4���4��S� �2�S�d;b_��~����q@��{ǔ���3�ko���Eh�ܓ:B�2��.��J���2�.��Ϲ_}����3���Ť�ܫ̇��r�\Щ�u����G��#�55�\5 �t�\{'���5#F��)�	�>D?�� y��Z{YO�m@FT�Lz
M��l0^Z��{lh�x����a�v]��~�o��R�k�v\�@�i��{��=1q���=t8�=}K�.UڱC�hnuN�[ӏP�����p�B,ݡ��k�����B��q�g���w�x��!��Q��M&]z!�	T]���ļ0^�;����*|��j�#{��G��y�F��L>� �K�+b3�U��n`����V��N5d�H�O��S���0�x����B�_59�u�D�����O_J*)<쮃��z�L��E��i$��@=%?�E��j�P�c1�bE�v�\�T��Ƭ�-ʬARzS[�Gje{���8��2.���g�w	/�rԣhW]�8�x' �����j�g��C65���e?ߥ�W�"�y�Q�|���R�q�6���kHS��I�.�j����;va��)Ũ���Y<�0%)#J�C��>h�/��K�nj�r���h�T�2"�-�"Pc�[B	&H�v�q$1Qa��a�A>RAZ��H�5�Zd؟��|�gѮ@7����GМ��y�Z/c?Be���3��F��s�(Y�To=�п��BgTy
��8��
����ȋhA��
A�;�~J5y�iG�97v��Oq��'���wAk|T��r(����X�`=�u#e#C���t�H p	}ѹU?�"��`Y1�w�+;
�Ue2�q�����:�c�~mzq��[����[��R����=���N5�K�������8d����r����fI����X0�Z�B��z��ץ�� ���b<Z�W��}�AUa�ȝ���lh�[Cw�b��*,�ń��X�Q�o#�.�b�VSIL��fE>*���ᢢ~y�ޒ]�7Ņ��|ID�id-e#{  �Bt�B@�.�����d�.k�!�2�I��םȞ�ְ�FV���ih�jD�?h��w󡋥|#.ö/L=I����L2�E�<��Ԓ�H��JԋS�MW��*n㨲p{SC��]m���-�աe&b.�_��暔ńdHz�0�����	���B}�Z����y�wOJw0�
�4aA�P_��SG`�@~��T?NO�i��yi�n�8h�d�5��%���d\3=*Xc�p�F�f����A�J$�m4ot!�:u����mK���y6�X@�o�V�|��n�#K�П&����Ĵlikn�Ę���N�#��{�G<��ѿ�2�D���.=M�H�(����ж�D����l��x���w�?&���Lp��#��M݄�5�|���l	�3��M�1��ɵ �Q��DMa|Y���ɊDivj��H@3�2~0���c���@Úx�E��yr'�r��̾�F7]�F��N-��ge!��0y��NA�!:�M��֕�2PaݘZ7��f0��ˍ"�������6k���G}��������qa]�z�򏥿.0���� ��c��}ZꙘ��^�@y�Aw�:�=�H�xʨ�V����m� F�B���j���P�R�M��wG�l��
����� ��_��X��UwZ�F;�p�8Aч�[�L��:���2b�'C�gӜץVX�
%�
hy�M�uE�K��	���=��F�:������n���<4�!�C�0�`͹(�d�kp0$�)wbi������j[]g;G�ϯn�-�_�4�o��&x� R#]��b1��}8!9�#Y��7:7]\�����R͍T�?�?y~u�ɡ,?��Q��41`?�&��W_����(��c��s����Q9+�x��M�'��GC�ԅ�� ���i_���Q�1�p�ggs	�E���I�ml�i���=��0�<^��>7���G����9�l�!}b�54�%L�]@09xB����;�������=t�P�#�T�u��[�e�U�{���z�?��:�qa�<�z�C�T��E�� gL^'�ʸp�cO�7�>Y��Yԇ��'R8u�p������L��=��M��>1�#��6IJ���>�Pi��l�'\B/�>����|'�ք��k=�E������ʣB�	asêp ����1P�	����n�>G��u� ���R���- �{���r��q�]"ǔ�N��G�#s&K�Ʒ�
�J��Lt�e>�)2R/7M��Äu�u���~��B�C�:9���' 9g���՟��%��8���h~ܰ�r������
:K��B�"
5c�Y��|��W�qe�F�0#�bKG��|zN��c�vS)� �@�f��Ԙ�h:֑�1$^�oJvHQ$��_�"�����X>��#"���������=�=��ڬe!�P�s[L_����;J�4������eŝ�9��<W	b�M����w~6�)^%�z+��G,�ӳ)�g�C�P7�T�D���0&��:�x���AGn�Q���a+��r��.R�g��N�;��`5)��_�/=� m<;�m*l�J�2`��w$J4B8�qܞsfd�c����B|��0�����ʆ&�̲i>x���H��J$D�#mH����f	b*��q����O�\���G�H��@��/WD��`�;�6�)�^e�0�0�Y�F*0��
9�h��$M�m0C��u���n���P	�72�Pd�ܣ���(����T��$w�*�o���Zx�ǩm�.rv����%nJn�%
���*~8��/Bɍf?4�	H���g]�dޒA8�<K����;�nܾ������#Uڲ+>�[�ڽ'�LPP����û��j���ȝ�g��IڻT���\6�M@��b�#��$�P& o�K�W���((Lr�`�l?ι��l�`�{�F���Ј�G&�<�Y��@��#G�y8�N2�a7(F�۸�`.!R����Z�B�E����K��p���	��C���FN3p{��m�r�%.�j4J�\W�ud�\��j�m�Gb�f
��i�:@��85 ���
I��K2}"!ՠ�2:�=$P_����V�!q�}�5xq>5{���
����������y�:�t��>k^ąU�"cjQw)�s�V���@n�JQ.�TJ?�B�`haDzT=��$j��kr�5��������eTkǲN�~�h�צ�?�J�d�����*�u6Oظu;�X�� �"���<���cj`]�l�qC%v��4 N��ӗ\�i�	�H��'÷X�Ua�Q �JJv��n �`����V�.������){��\�8���O�u#��Y��bM�J�CO��Ν�u3���� �(�h��\xVSAv �?����j��&��)�ُ!�\�э:
�X<��B|�A���u{���n�������@���Q�w�	nb��� ����PI��&�/���$�J!L����T?;��sل��$(.�a�=������h�+�N@w��%>)e����U��<��߷�(T���nN�dN-��crj^v�!�	�����/fS]Ȣ΅��Zu0���	�b�Z b`1�![A�o��m�J62>e����{yd~�8��$݂I�Q��GC��}�G�K��p�g��G�/|sM�D����{��K�����^-�%��?3TgFz&�Pkgj-K�R� W���KI�5n�c���
�����gC4��A��_7�OK�ؤ�D����	�0SSwO�ɓ�����VP�z��������MK�e�87�I�L�VV��P���XKz;�K$f��eF����A���@�	��ن���e�֞�x>&��2��K� ��|���^���\���Q���SD��a )�.�%%���?7�rG�E�˺Vm"�=����:�X��j�5�b��]K��'�xOO��S���e��j��@����!���\ڨ㊨� I@�(+�����3���OY�Q���</� �X��k��=�Z�_S�ϐ�����oQ����&�U�;��.O&d��f����P�>�BNEi׼�#J� A�����
9 Al3H~��wng�`BS�q�J7wW2&��i[a$��mS��o���>[I�O��V��W�1WRlY�$�������0�o��^�E&�L���Y��qCӎT���N6gTn�^_�qM�9[�aW{�&����8���y�(��8o6I��-fm��kh��QLX넍@��W�%lכ���!�ϣ�s���tq(�DY����J��{�>���l=68�9��!��T4
r�Psr��"��]ï�lR	A�o�����H�|{~3�X� C�C{j-��CJ��!P��D��}���˧ܝ�8bF.����Ԟ��f�R%|�4n-���q{ko4)4���T�ԃ��E�
�S�Ţ�~�T �@��U��He�[;d��&�9n�����U_�5^��
���7*v曈��b��<3�V�,Y��{ZM�q� ��6x��.9׿q�{^����P����D`<Z#�D���TY@ء��%B��T
�r*{�4.��b菸����B�ӊ�pI�7�?Y�b3>�#o�.�u��'�#F�����*
�t9͕�`+ڙ�Z���2�7)��[^5Ÿ��~j���ՆaE$�(@{��|���(����#�������L���P���ǂd��bCs3nń�~ae�b
C@E3'�P#5湶�ǣWȷ�Խ�M?�c�� ��s5@�/�2�z���H������CL���&M�S_�G ���}�ӛ��L�ͣ>�����u�V�ud�#���4E�����z��E�ױ8Q�������+0�=o#J�zm��<���L�6��4��Y�s������pF�C�@�V�jd�rm���L�(g?z.o�E���v�sQL��Q�:S�@��ǁ��Қ�#��i?���O���c!
��}�:�����LNY��d �n�����1D��h	ʰdd�xn������+�7R.���&��(�M�
�p�kwV����7���W���C��|\�0��CRX`�< '���,%ڢd��T�^��!E����]��]��Qt�WKc��֐�Pf�U��g���7��$��\�1a�)v7�k��-"�U��8��*�-�^ׯLˠ���v��$QO�O��;�����O�R�;��Q~:�a%uo�R�PG���:u
��;�?����9T]f�C����:��㗼8�E��119�~��}�n�j"eӷ�� ��h�R=����[�����L�}:AΌ�6��|�(���be�lG_𧍸Z�ș��UD�����7�Inrf�9�����6h��_��b��e�����+�\���)X�@�|d���e�\ ��x2�����p)�q����z��~QE
��![g�����H�9�]�e�$L�m��)�'�_��F[Q�7�
�v��L��e��S�M�3h����dV�`��xm�OŨ4EC_�Fa}f,��^88�Cw�թ�ts\��;_��l �8�H��쯾	[�/�?46�,�]y�䖩����`�ǹ�C�M�L/���E��y�Q��m���Զ�9�V�_1���������&)v%�+֢mzeK,s	����5T*���y�=�i���rm�h�O�h�v�8 _�``P��f����q��9Ý�S�y�dh��'��(nH��E^`�RU��j&�8�v|)�q�D������^VeY�R\�U�3����a�tF��@؋<�ԃ��E����-r���dj���� y�!_'����'�+3?ꓸOצ�<���[�؍ &g��F��������ǐq��+�1$����au��5[��@��FY<<�]a>�n��.�/����v�.�^.9�%��Q���PT2G�.�*@v.�؏{o����=K:i�N�b_���>:omXb�Gb_��t���D9�Ms�� ����5ڵ��M�۷puf ��e �>Yܵ��9�R�7bů���r�)�B�5aaR�ڥ�����uxEN�sz��%kl*��0�`�u����@1���ϵ_����0��_E��"�f=�r�#��j�6A7apf%2�|b�d�d�۟GG�!CwY)K�0��~��XQ�U���[WÅ��� x1`
�_��Y7*�fD]��
�����DV��޶&���5{%�U1�1f����u����S໴<��x�IC<�%�E�dIv��ne�VF���m�����L�/�~łwj�'*�WT�_B���t�rr�$O^WڕlL�/����ڠ��"��8��۩9-P�3��6w{��p�8�����T_���c�qy�2�~�O�9���:|�}=U8�=�W�y���25�k��2�sJØh$S'yQ�r7_��ǱS<G�h��6q��X��b�h�h�jL�|XRz�?���-��'Em�C�6~��46�;��,`����mЋP*��H:ﺼWrt+�¦x�lJ0�ݎ�'+��������='��n]�;�e5G�B��ԇւti����"K�ŵ�L����b� oe�*�7�10;y%��+�zI~��BF�b6m� }0��/�/�T��^�r�42P{ ٦� ���ό���H���՛E��4��:2�%����Y���Q����q�v&��7�6�Ģa`��N�غ���:�;H�D����a���Nal��t��#��V,�Ї)y$%�Ҁ�䮝������xGU���:�u���
ʀc��w��|�@g/��w�����Zi��NN�9I!�݉��cI��&�ݔqv���F��ձ�di�X��Ah��'�� ����\ς�嬅�rJ���lœ��ŬD�:O�{!{�
#�o�Ѿa�����j�0V���ͯ63�-�Į0g��TI��S�q?!����|y<��6�$��s��l銵!�^�Y��\��AV>n�{P� (�[־�%6`�Ǻq�s����Ċ{�"~�,�	�t��?�I���/�f^ZN���"���q����U~�7����Y]�b>�B�xm�u�ľ|]�1��Ոؓ^�U��-h������ �n�Vu�O�ꕫ�*mh2��+��a�	�N�� ��Ҭ�q�, �팶XM�4�k�]Eԡ�a�	`�q��Ĝ˴�	4up�'�oW����6S�(�	o�W��! }9>ަ��?{�B�|բ$T )�������%ا�OUm'�����%�du������M_�9��ue�u�|���z7W3)?�d��k:r+Y�n�������(5�k�>����#�J��-j�fs`&�`�� u[��`4򯉘��l��/��},�ϖ�I�����!(�,�m
�]�F�Y�%�G�o�mqݝr#�af4�i"��)�:�u����Ni��m}�yͫ́��Z�! ����ԗ��y	ؼ��B������ϔt�P[�_ݭ6��b�d�EMt��e�Dn���V���,ד4��BH!��(��#ތg>
����}�4��.,��kU��R�I���~����s.w�h;�v�r�o>3�l�	��� Ұ��B0B�ϼI�Z��0O�~�_���3��t�/MyE�CV����7�iͩW����=Н��ِl�x�p]3wh���.,�U�lJD��8r�yH�G��Jç%(�{'K�]@�x	�x�V���wv��I	=/ Bb�!x@���AY|���f���=��BD>#+H�Z{2���&;)E'��]����ly�D3ldwq�H� ��S����/�7Qަ>�{�1Cd7)Ev�L���l8�����)u��xqU)�1�<�λ�?R�Vz�S��S��z��-^��cjl�X�F9o�Zx`�1Q��YN$Z�葬r�
/oe���H6�=����^�9ѝ�L�Zb����A��]�9o�M�b��L,&��� ��p����,�l�e�;}
�IJm;�F��Y�4����׬~�Ư7��'��y��I�9���t�h`����XOyڮg��a3��\ŋ������+��,`h����ͮ	��;�r�j�T#�ӷ�&��N�Q���;�`aF�u��A�(^�6R[}zm��U��(딹��8��,m>��bTF�$��뻿׻�I��Ǻ��e�Q��/�$'@��/�ɬs��	���$���eP��?A�3��O��z�yڑ�M����<[��՜*��0%��e�9���CgN��y[��	��[��E���9k���$���f@GH?K�%zz���x}K�}]� g�}D����L�� �e�(n�u�:I�O��9�����W E�dF�'_�잨�@����	 {��\+��z�bO�����;w ��������'���LU�Ą�V�Bb�ܞ׻B~������\3��뫅^��u����,����+x��o\�ֺC�&�}j�4Ɛbe���:"a�W�'�5�O�џC$�ޱz5������DYJ_�&shn���	�.�Ax��WW����A���z��Dw����h���F	-W��]�6��}�1�Lc�����V9N6�^�>�C~	k�Pљt�zø�<��u�''��R����hɨ<�`�Ը�m[X.�!���4b#K��R��5:O�7?��f�=���|�򎌟;�ä��S6N=��6i<."/�6����㼛��S�o� �̠[z1�Q#缄�_]9d�H0�՝�h�R�t����gB� r;U�v�Hm�� N/�z��r����|�O�����i��_��}rHEZ��VYw�Q�Р����a�}��ZoaX�����>��@�\n��l������zI'�_���]o�},Y�l�+��3���!5��6w�����M[ Z
�? �g�����}�;�_t���Ɨj�"�@�jX���#JЋ��|ڱl|k���i�햋1�Ҭ�nVL|d��?���_��W8c�+�uxԌ�	$�\&Q�z�����:Z�E�d�����(�� ��D��vZ�,(d���S�q��ݕ{h�D!��-Y��g	�t�L�F%���ԥ3b曀���w�EBa0RH�-���h����Rb�
���X������K(��$� Y�97�Q��FҘ	O�q�����9��K
�7X��S�8�(g�&��{�����Q? L)�y����qJg;�b|�VG�G��扎;��ڎ��̟>���~���I z2x��Q�)�ZP�l�N�P�~���PC�g%#����
��Y��e������9�(y��Gd���� p�MX�������4�	,ѭ�NMʐ/�i�ī	t`�R�vu��i�@�Y��[j9ijQo����@��KX�f��.�X�!zu����[��nVaIt]O>�C�=��N�hG�K���kES���0��6}jrPʚ��7y��Gp&lm��Wiӣ����+���u�x֤�}N��Uc>�\1�E"���;��F�\�������zv�s,�cH���A��{�x��|L0m���Zy��_3�����twwQ�Y\jf��+�����ب�%^ ��ӏ~6���k����1dV	�����ГB��0㠴�Y� �P{`�Nԝ7�Gw+ȿ9W��������ge�?,��׎B��L����g�zoy�|`�������Q�{bݿ���д?���j9��q�B�$����D[�Y{����6�9�?X_�I/P�`�o}>�P$����D}�������D��P�4#�!�	��gQ�{J/կa�e�ܣxoA�v��\��K0�9p��Db6���t�0�=��˘M��h)%sҥ]_���̧}_�!�F�h039D���aJ�Ea�1Q��b`��Vb��7YGPO���I�^�uY��<�PF8BAϱW� 	��0u��.�ɐls&$���[��V�ΰ�>FG#��2��D���G����P6��63�*R�]O2$���>k���q&"��w%l߆�Jƫ����^��cV0��@���)�pRr(~���<�91��:�\H�|��eMTk�EL��^E��y'5h���s^@m� ��O>AR��cF[O���-Ņ����cs��pW�Ù/-�������"�Khk~�� К+~6��m��e���h������޵�O�YJ{��e�Jqd&h^�]��<63��U��ݼ�po�M(��!��k��6ç�q�,��0Þܞ��j��&t�a�����1	_���-k�k�w���=q�,�i�X�q�"�u{�}�p�Q!ǒ�ܼ�y�QX�$�/����}�̡F�L��Z#��cߣK�	q�T�و��!���/B�C\�t۔�j�&{Z�qZyj���&%B�pY�]���vR;ѕ��D�ȓon������'p�fƱ����h�):o����IB��������r�*�������Qb�0�d�7(�xws��FÓl�<�V��fC,�G��	��8�V2�r�̒�
��A��737��#��2�&�.+C����%�	50�����rN��Ȝ�1����R/���)@	.�Zħ{�����P��(H t�R��k�;�LC��w^���|�/E�\��)��C������#,��"��o�C�q����(Rcb��`�3����[X�]��� M�b�*�l�&�g�0��K����جFD��=u�U��"&j��v��t^no.n���b�<��=�W��'��~�r���"�	���+���!V�$��3��Y[Y��&�������L;c6��{:��eQ�$��,rsH�\S� I�h�f���V��z�F�0���=(_b�Fv�\��{;a��Ht�tbWnOP\��U�L��d��(ᾱ��S�����si� �|���*@�w�P"mf@#�ƭ.��g��B�Q����(\��M��>H�-�{"uFɟ����T�Y`dg�vt���f^.3�}��y��
֧��"��pܓ��k�����J�EV�P��j�<��&���?%P �^�t�ݿԲ$��2��G7p�;��SK�Ia����JP"�2X�'=�����{��F���鷆���zw^�v%T�H��6ӠҦC�[�m0-ȍ,��/	u,�;X�?��+@��3���g�����Y-����3�㪷-0t��Rg
�J����ש�ԚV@ ���Ų-n�^�GQ��E"7������!R�>9��#o�&��ю呋�F2t�f����<J�H�0l�$�R�z�#���iDJ.�"5D34��/��b�V���V��B}C��;#�0��~l��Ė�?A�-s9���$|ͨ�]�i�+6��TF9���(���gs�����G��C���C{T�nV�� S��V��T������U�TH�����&#ˢ�A�ЍVן
������V�����yp�lX?��S�u�5jG��tOh5%�m�J���,�k��xR�a�H��#+��4@[�����ZQD�&��SY=����o��ם�^-F˻�8ep������"���H�r�;��󟀋�v&�晚↗���h�@1!�qӮ����oV%J!�t3􊏽�7�C7���G�=y>���n�Ʋݽ(��d�	"�n?X1��sk�(jѹ,<��'Ό�wc&��ʣ˧�T���q�iM��B�iqA��</���O~�,�T��hN1���2�%E:}<����e��P�J�������_�b�[���q�,�}�ߧFe��ʫmUd�&X������>�BpYhH~�L�dլg�#Et/M�Vs�O8כB󽜚1E���"G��6����d���%��F��}�Cט�{��Ľ9.�Q.4A��a��&�5�M�kJ�I�)��Y_N^R.4R�[٥S�a	^� ICEBE(���j춝K��&�7�����O��t>N����5����K:��O�`��j��~%�Pƻa��*{f���͛��BQE~�7 øy�o����nE]��A�P+���)�V��~�r�a�*�ꖗ!{�� KaY����3A���;�,ݿ���W ����HfOr�f�p��7g$( \�Y2a��r� gɟ�[�J�?a^�B	"��9c8�5|�A�&Qn��|gOi�>��Ԫ�R�y�q�y�S���$���P|�����4,8�ξ�,EB<���X�#K�0����C
;G7�h]�;>�ی�n]�S�Woo5��+1�Cn��K��0˹���U9���n,W�&ه��MK0[���z���]J���9o�~��ܚF6uKy�&��a�=b'zd_�e����Һ@og'P�a�$��P�����mLc(EM����$M��ȶ�S,t��>Z1Ř&�͝M7PnZ9L+>/!��I#��|$5N�U���Pjcf���D[��;[�gO�:/ZC��?oA�ȏ�2�`*�o8u9,�Ӯ)�'��F����&� �66��6&���ι���uwREQ\`&��|T�g�K�-O�t1�#w$w�C3�T��S��&�B#˼����"2�K�YG�{����6*��1B2����h�A�@됦g�͚�����[�`�'��^�͘yFK�Z�WD�n׸�79m�0�覄%��+����-���o��8ũ'u�YM����D4�u�yi�H������^����(����R]=�9���]{+&��*�"�3\0� ��.���jRQ�I�+B�F��.;%�뿨&��	����K3����>�M k�3��F� <)0[��7�7���Z;�ظt��ݥ ��~�(��~��kI'��(9Ѥ��UJTr�vk<�i%@.�Z�3�y,����ϊ?�7L�)(���ķ���}��+`P���}���7{ES�ׯܰt;��G���A8�Y���^VnU�":�����Hɪq��F�������1��W��TKkJ��t�}O�`eXJ����	�]i<�&�������ڷA�ڞ����(�;��
���a�n�x��c3rK�[%&��cI3+�Tɷ�7�H�%/�p�ֱ�m��|H���
��n�
�z
xwy�H�?CTD��d�>6�2߫�c�OK�yJ@�ʅ�y�ǛU3@-he|�|�@����B��7j�A����}V�^��G��Ks�L`vt�Qa��|�����ycCo2`��qYJL�Y�L�~�Y𿗀�)R��3ǰ�:��_X4�Q�c�&��^�
�#�t�q���F>�I;� Vd��h�pA��S'��9ѕ>ZD\͒��,��k��+OhG��5��� �ѮK�<P�hF�!.��ogn��r.R]Ra�a2�<x30�N~p۩������B�u)�H��D岵� ���lJ!!!Wv{�����ј����v�z�,���	��H+�/����n2,]��@X�!m��5�7��w���o1�V6�W��r�ɜ$���� ��}�ix�Y�&#���f��~��:�e?����x%��ZH]��yr5�4�<��X=Y`h,d�D^z�5K���%�Hdu@Ph�����Ľ�ú0�W�����k�k�g�}GJ|�?JOb
��)zЧ��O 5w�}��Bc?z����Z���\�S�f�g-� �J���Nft�W�rC�1~�C��(�?�Z.hq��1+EҧR��G��?� ��M��3b�/�9�J���lЙ������%?╲�`���ö��&y��t"���؂� ��jv�C����ً�� u���Rn��oĽv�D[�� \u�G�AĚ�b�J����#�EV��Y0�ܾ��#�z<���x����y���J�$힅R�P% x�������QT�:4��jљF��W�̌!Z�mEAʢס1���`A[5�i���q%�핆��1�靜��¨s����^y"��u��x̧ݡ��$��i���������V��Aw��<8��S'���4�c�4�A˅�����F/s#�M�ԣ��s]�CU���j��f��\�����|�9��
E�8ʣ^�z�SgM�����]��.��/{J��G�
׹e����_<�/�7�G}��1���V5x�hq;�����Y㇏��+eL�Sb�z�j=���n�E��ZAR|
q-��C6�Hz�u��q���e�#8�R����Ɯb>):0�N�����jc��O��2��H��ןi'�8҃B��T��{P]I�lj�q��v���乗yK{�3�6�+�8��)�	���s�v�?�TN�ŀj̡S(�R����NA�Z~�
��-���"�z�!�x����ȅ���rx�B�0٤�g%$tN�Do7���+	���m#��DE�\H�wg���J�M�NN�!"��c.�+�A'S7�9���Ǭ���Ι�)ʏ��z[V3R������S%�����$�?�A����aÂ�Y���S�P����`7.wo.��2/XHo?�u���Ǿ`����`�(-|�	���ӓ�@CcZ�����n�z�GU���n�zN�h��-��,��2{��O1����g��H'�B	��-C�Q��ʉ��)�{�c���.�h$"�����aw��-E3B1J)�����s�C�°^ ��(�~��Hd)
��CzS�ջ�%U ��XHh�A��a����e���/dJ�H
w�
Y."5C�:�X����(k�����t"�}��wl�����9�*[�0�]ꭵ�R :�Ժ�v���*�_��a9䝠1�����@��:���^�Ԑ{���=-�	W��U��p[��=�(�X{��˳�.� �s�)�M;�Q��X��(Ø�Q�aJt*LIL/��{<�jT���j��u�_��h"�{�E���+n��L������?l��Q<Ϣ����j����n�k25ċ��gv���K7Bۀp�u�'"fx&�.j[a8bu�{&�}5�Z�<A���5Tc�z�-�
Kn��$f�*^��jZ����Y��xZ�g'j���0���$s��]�$֓�є魱vG-�z�G��:�iVT׫��-���*\���	?�nSżv����k��R�V�z�DS0�t�/cV�9��R�V�Br�f�I��\���g��е�pۥ�Sw�s{L�,r��ڭ����>�j���}N~'�(�Fy: pƯ�`*��zn4�W��4)�*�Kx���XA��X�AȮ�<�5���&)}q*D����W��٦|W�*�q�`�s��X�_yY��Ďz�����[芣T�C҉�U!9�;���ͳ��2eZ�'~d�����t�|�'��t/'X�sknH�@���L�U4<�0�q/�&e��e e�q��X1���^YCj%�p���/i<G�'��\��,`�E��s�1����nF�ێ�����$k��zlnT���Dj�D�2�UMuۆ�}B���*Ѥ�E�:�O#���EQf�P��".�E :1�W�Z5��ſbѸ�"-#؝�?H����?�;EYl��tιSv6�n��[�߂V��˛Τ����HRJan�ɦ���"��_��@
���PWq��~�[������q��N�h.�1�dB>�Y-�c�'E��[W߬�Q�/��� ��L)C����Ȩ�<9�;����m(�=}�&r����?�&S���Ok����z�p��X;%��}m/VQz�s1�ip��x��t{]��K؃��@����+'��K��p�PXgx�O/@?��{cB�_��f���Lu�N��g��s������¹~���eֿ����4�7�2!1���lHp������^c�7C� ��L����G}-4��݂�@��v�i�v��G<��,_Ls3�Ѕ%�[@ K��U� �d%&��M�<P�Z�J=N�a��U�/�0�����E�]@I�CGJ
��s�1I�[i�%�4��!,��r!�A���|�,!�g:�Sb���Yo寬�E5M***6;�>�6�5Kxs,�nn}���������� ȇ����֌]�������_��5��<��j�1Ց�-=��W����{���0"��I�Mr$���Mjp�n%����q��p���blpЉ��+��'�X^���u�C��JuH'C�S։^�=u5�:g	xI����}n?|��FK��Z6<��f�|���+)uQw$�������*`D@b�?w7�қV���@;��L� NjM�I YNW��	������9c�({��3x�@�A4d�:��e���/��癸�O������{+j�M$լ�UG��N��O���L�u����صFu��	��94 �v�ГxV�J�j���6d&sI���fS�N
z��j�6-��l�ͥru7�w�N��-KyM��eS��O��7,��l�U'��>~�>'��#��a��L����ô
������n�s�žY���En_��l^8ƦI2���G,������rz��;5���C� B �+�M�E�`ك�mg����>�;<��J�ν��>�T$C���e�=�⯾���&�����|ſ�u��K}`���_�\',~\="1�� o}�xAV#���ovtz����|��v��6򫍘������4�vݖ����0�z�,���L�=O�$��^����Ue��0ٚ� ����suxe#������=�U{ۡ_��ޓ{F r�e�jsR�'�6��p�Ct���me����'*�ub���'�A�a�� �֙9�P�M�1t��P��U*J)Z������Nݝ���?	�7lzC����H�S�]R��<�S�vV
BE0�S�5���n++�hC��e5�}�D������P��s�'�r���đU�9��W������#�n2�Xͣ����b=��AD3�s�Q0���������
�J6���1j�77kjz� ��������$C��X��2L�9��U&r1*��*�B-�R֝�����|����F����7���j.n��t����J��r��ۘ|n'�AH T?�j"R�N��6�%���mh�6 �����U`�Ό]u|��Il$#]m{l�Sc����^h�-8��8�c�K���y�F��a�&^M	��K��*�FV�u�|Z�>���P�S��v�?`.	A1��z�]�ñGjo��tZ�|��)��b��74��b��ܯ=r�+�f�6�)��m��X\�s	��yw�4(��,���O�Z���u��梨��\���7������5�E�*:*����SZ�r�����cS+\����(�	�=��q��S{!3�@d]��]����y�AYz�xl�Jp�%���k�i�2y5��kL|���Tz�4�\����W����(�SQ+�� �Q���jV���db6��g��`�Ga���JW�(s���`� 	��k�m8m�E|,��t��.Ro3FθfbTG��*�h�J<C5'����6�F٢�s�`���q���[��cl:�lk���Js��֙ �f��R%!&Cdߛ?CMe����i�p5�dw�r�#�zq��{n�'���֣��u\��f{���AwC牞]�xËJ���d*p 盦�tZoH�2-�{�wv�ܒ���J7�5H�p�e�&c��ٕ�路̅8k�x�2!�^��u���\�s�JYjP�J�1k�C����
�m�f��+���A1�/�Z"K½���ug��G���Dς�DH�Sǌ�{�g���i8���Ķw���}m��|h<I@�qj򙪅����b	&�DOZ�M�̗�"3��k�$�52�=!��ɢj�@�4��]�u��zfmpo���E�/,� �\#��(�Du��Wuӗ��+�4�qhYFw�t�<O��e�hҽ{iS�҄D�AD�_y�{�E#K�Scѥ�5w�ɾ��ʒ`9���W��>��Q����<7ݧ*�'��(��$�dJ��kqn�ޝ3뵒��W>P~4��H>�X�A\�����΅6���u�����yol9�
}���Gˎ~�v�z��+J��X!�Z�į�a��*�����_��k\���6�$��уs�:�^�0����K��]EIh�q��Fe���5��ў��� T@���F��ĭ�E;kb�ҳv������U���,����L����[�0�	�ӳrq��F|�,�]�%��8���n��TɈB�.�����Y-'�1Xw��{.�����qT?�+�8���x����4G#�|�}.��U&L�5 �yи��*؝�>��{$���&����{�4^e�G�l�84|`S��P�ٯ�D-�����՘R:�9T�O})�d-�9ru�k߮�����������lMƗ�O��Ŏ����&D**��"���S'u�zP�_�}$(~1��1�hG���[��r��ST���a˝x.�>V� 蚊vC��$�LЪ���5�5Y�&��+͌3~�.��s N,J�h��K�5-�h�Pm�g�e�?��&l-\8�B�����K�<s��H��hd�m�|��D��qo=�\�z
7 <	:;��Q][�n~�X��m������ej�<�.��$Z�� ~�E7.&��Ǎm�<b,F�;e�SX3��m�FY�JG�T��}��'���g���Q�y����1�<8�/	7�Qq��TE%Y��{?��.Y)d�y�&���.R�x�"��GN#��%�Ter��	(\/�?7���;�}��A��v66�k���c�P+M�do1Gd��H�p�� +�}�d�"z�&�;cR�&�ܶ�CE�ڿ?&͜y�Yޘd���/Rs�����+�9sc[���RG&�0h��(�3~M�F�9@�n�*#���B��v8��C�ѽ�e��E�Ð���z�p�Ey��ѡ�U�>/�%k�/����蝌�Ŀ0)H؇_�ř�0Q��@pV���O�°r����ˈ��p�VI�%Ҍ��v	Y�w�4͏�
���l�/�j{�	��
a٨�GM3v���CI���O�!l7ׄ��)o���G�'�}�ong/e'����r��h@��
VĽ���2$�n�-pl��<�uWћW_q�7��>R�Ɠ��j�1�UC4�6���z#&M�_�wO�]5�~�˾j��
k���:��'���m>ܓ���tI0�1���%���Z��0ͱv��N~]&�����Y��^7�(RV��	��_��r��If/a]7���O?�@�{fx�Qb�w�F�.�W��<1��Cl~�
�G�4����W�K�'�N�҃��=����W�(���`�G<9�PpW�Ǖ��ª;Q��*�������4XT-.1 >���?�,�1�
T��G7'�]�c�v�׀6p�8����m�\��[�
rÍ�g$y7���s�x�1�
_l���D�� �>פf�s<�Ix�t�hDx՘s&Y���v� ܷRr��[��w��K*����i��z�,��Q���}Cz1/�+:��ѩ ~����9���I�z�#��J���e��_�b�I�$St��CC༁�I�tO���#|w'��f����>�y(�7�X��757~�,�9Z��}�A�7f��,��m��Hj��&+�
p��V�F�)�0b1�D z"���*خ�J��gw$�n�S�b-ր�kP���>kl�pS��e���!; �9�j�W�����^4ڹp�éќ36����p��������[u�����y`VEf{�>aW�i�	ȱ���YE�!�)E�/�!�VU0��iu�^���sȳi�� n%n}�}W�4h���ԃ�*Mb4AS��1�q 	��J�����r�r�֬�� *���K��'��؎I�r0��l)E�=	}M���`)���g���&���,��jLN�W���l�����-�=��r��X`f�L\}��ǂ�<6Woͻ��P��R6���^�f�-�w��9�)�[�����	���Vƌ�Z}M��t]�0D�H0�W�,\8^/�H77�d�TE�qsH���F���U���LږR4�[�o����^�E��::�{�;�'�0k`G��X
�>}(�a{5|���B�<O�xUׅ ?ͣ��)����A�-��KQ��'h�&����" ,�(���Ä$�%���i�yn��'���Ɉb��{)bX�_׵t�@|�<Ҩ�4�EޗE�u���l����&���r����W�IZ�F�&_�R�8f<�9�h2!���T1������U�l��Y�o6d2�*��\�F$+Q�#Xb��m�#y?Nc��rq1�F-�%fEj5
q�$��@I����� ��~�&�D�IW��˻*rƁ3��D����� ;��� R�|�,g�3����5�q�YZ�6�����N���(�xU&�`,>;!�R��j��%�w�v��GL�/^���5�a�j���4�2��zp	��E�[���C�t��!s����O�1/��.����'��o�����<�`'_�z����X�qQ
�z2�0a�/�d��Ь�ap]�Y�9��k� �e����(W���2�kڪb���,U0�8��~k�xz�׃�w��bw�8l�BO�{0�I;# �lA	�����b�nZ'��`#X���H�3Ca���7//Md\s���P�aP�h��|���qG�D��C`�F���g�i����Р"���.�"�=�� �\�0����qK���ސ$��t�M����X���3i� @�ԡhfIm�A<�ӹ ��,N���=�v���+��t@=I�nk<�ǣ��i��WȮ��E�k��	����]��֫Kn�jsz�I�����y�"���t�oU�x�y$9x�n_�N^�=���I)���*E��h�}#г��T���I�m�z��u�e�����=KCy�|s��V�]K?��X�錓W"���[��V=z�<WA�}�b�h6-5�}vPsP�+.��Rl������6E���w��W�t�~��n�&�y�"х?�*�fP6Yc��A�S�8:���J�4(B��dh�^�ٌ��u��L����c�CP�T�kM&R�+ċ.U�v�k��E�t�:�)N,�ǲ�"��|�ª�E'�)���OL@���[�$c6��q�7/K&5ɋ,�?է\H92�l��Z�pT��S0�(�ss�%��Ӣ��7*��D�J�S�MB�����r{+E�no�� v���P;�gy2��@�>O��:KQ� U�7�9�;���.�b,h않?7�f���|���7Ґ.���
\D�t�y��X]=�����J�*BL�?�>�>����7!z�(��K�S�`�(2
�J���� �*����炞k,�`�J����f�=.���ݦաӀ�gŐG\P������	��\�Q��[Բ&�yQ?7�Ľ1��l��ެN�+uQ|a��Gg����E#V��5]�o	r�m_����x��oC��2���<�5��^v�07z��[��n�c�:��XY��K̂��TS�d��N�i
�܃by�P�.[����ՠ���V$��
�V�v���'2���Paw�r����l�S!�.4)dҞݑ��{�����@��~���r���:���Ȓ�B��:JrA�n�����(��O����<��R�q��I����a�O�rn���)!k�r��%���/╬�2��5������&^�0����2��>"N��cF��1p�yJP�J2�?$�(��}}Rap�1��d�xt�'�U��֔�͊p���u�}�����]�pF�h��*LS""�/��5h�GF��;��@ƙ�������E���k5��S]�yU��uFJZ��m�b/q�+�tN/��V	G�?ǥu^\aC�h�73�WS=.�:�Kw"��%�V:��1����u�)|��?�n���%%,M���u�gAn��y�N4����*dSN�&1diyi�1\U��SO�Q�K�{�-w���;U3���8�;L3ATb.�ٔ���O�
+��Q��i��կTn�K[ɑ��O/�q���M�ُY�_�m�����Jbs�Nּ2����ΛYFIi�
�[@501�}�m����K�����库��w���\�(��+���ώ�����J����h�#2��>V���,�S��
�o�R[��K��U���,	�T#􍼩|y�R�.CBγ3��7ҍh)�0��{�~�kUr��g*N�Ua����hX-���-{(qF�O����V�CH!@�+=)#�#�]tl�V����!!�\2��z��xk��]�h�$�\ؐ3�1}Ё=���/er29�
�b%��퐡 4eh���ڑEd>�h����n`w@Q:�ՙ�9�١XOy�GD��G؋�RLy��2���<��ok�.�S����YM��4*�iZu*��7�9S�"l~5/��9TA�ޭ`�V���ƾX9`�<[��˄|}����/��8�l��;b�i�F5y�'��W|8^�L��<@���K��K���ߤ���K~g0��7f����Ft`	��MRً�]CLcd�uL�ॳ\m�*�5���e���_�p��_to���1)�D��˴�ˀ-�3�|��&^M�h�)�k��^?Vy��d�ZQ�����mj�e����@VW��q{��sxҢ�~�.�^_�܂B~���
xFj� _I�.��|��A��H��c�յ�YV���,���h�q�fp��X,�aVݛ�/�'�0m��fV�}���6{A��B)��wkT�����amb�B��_�YI�<Z�7�g�ܼLF_vHZ����JR����`�	O<�>iu"z�J�(��y:[X[
j����D�r�kf,sk��$3�qio����#:<��c�s��A�C�����]�B�L�'�u+7M�,��}�C,4)����J.��ȉ��4#�^����1Sh%��d�����9Ʈ:O]�����t��UoE�	2�
��`dhq��t�wg�N��R��Z�w�K\���D��UQyV>fC���_�$1%��ԕW�ц���k����N���(4A7�W��g�i�Iʆq�мj��F�t('�OH�,9�Y�2��B�'H'����9gA�jA3�7�E�����W��,=sS0����y�dDY��TF{7I�|f����D[0![{0AKk���q����2���A&�}�^����4N���w�ش`�f�`)�n�Z��b��D�U6Q���㣡h��AU,��F��Ύdhh�$]^�����a��6�R������q��|k'�Ue��.�����a�U���6��R~X�-ib�I/�����n�(���;�H3	����bu��)5d%ϡ}L�,B#�\��K�¤v<T�(�� �-Nǔ,	+n	��N;�R�h�����ZH#鄫S��N_��EF�嚵r�Lw�[{�N Ԭ�T0t�NG��#�������@6�(
:~l-�?[�E;L�/8Y�E����G�p�/�@o{����)3�����?�ܻt�3���Z�{�L)�"�>�Ct�}3ja���r����d��k�ք�ux��pv�EGk�l:�a���b�;�"��83@�|���a�Ǐ*�a�U�X6*��u ���,t�Jb���=�o�$榈�dD��>���+�&��[���4߁w�g���K���
1ˮ;�� ��eu& P7YV��a�?@n����"�˹��C��Z�T;�.!N��	}�YZ�B�#�NC@���^Z�R(]rV�ޠONO��z#>�Ij���~r+c
[���ƽ)���$��-��NJ1�y_�b�,Xن��{��38��,�1�p9kk�Ai1H�q;��}�렩��j��R��&tp�J� V�B���# �nY�1� �>9�Թ�pz���Ԟ���ϋ3�W�]��Bc�-:�0�Eh�mAj(;>?�����_��"����i����&�	Q$6��`�3>Q)�agC��iQ�L^M� <�h���k������9܌>S��,f�zk�4.�h���;N���P}�LM>yT�Ai�Y��L@�l
}���6�\*����h/-,Rp�C�]����O>�ꗵv���x�Q�l���a�V�pD�x�
J��=ߦ"vԅb�M��� ¿p�e�䢵l����8�I�N�K�sҳ��_�����^X�w�md���[V��;l���f�g�8��gc�Pia�X���ߗp�5s�s��*iL{Pw$P�L�ڡ2v���T^��P���	� �F���dʳBR��%�X��QY3���F�b@�0�C�D������	�K��Gj= Bbq��/R���q�*�B���ڭ�_��˒���RT���JD@0���l�{������K՟�,� +��p0Q��8E�i_��}��?+�'
��e��&�B�6��)ȯ�W�ǋN�ܯ�x��%
P�
,/�(h�1�8�b��A��K4���p�� c��5k�e�n�D�(��4m(�
��a���F�F�Pd����$H����)��P�6�vӑ|�c�ɯz隔�5p�l�_9^N1�r1c�06��4Nz�,�-U��*�$��"帶��@QfcFX�%[��r�$"Je��P�V�cE���P>T�JW��]�_��1r�隷M
L"�+�@���ORڝF�k���2���6lJo�z��S��[���(f�k.�e�މ���Cz)ɼn�k��fP.�5�K�W���E�k�+�d��tH�N7�D��Y+�:�g�S%u_`/�;ip��Ģ˃���K���L
2'��ōaW�PdN�����5�B�g1}3ҁ/I��*��1�4�fEC���}s�\?j9T�˔�BIU�K����]�������a�_���M��E�g#Mm<�%�q���fX�}��	���
�<@�f7���~t�<4d3���PH���?Y^��bxƊ�\(+Y�ǅ�@27�b%v�f~��{@�h\�Z�	��MK ^wk���]c[�e�Z���	����!x���yC2���:���wZ�>U�������[�����JC��0�MЙ]��zt��al����F>���ԣp ��E�����?�8����m�����wF C�5�L2z���}��y=��Uk��@U�Е"��N��[<�G��UJ<:H/��Π�W5�mYƢ����&{?w	Y�_4��e��;6nBv\F��/_̷3C9dh���g�����>�T�Kd\��#M�Ne%ͭ�.<����
|2Xٷ�c�6u��-ܧ���lm��;�o���'��K�0�$�IHm�����9dd]�V��Ȭ�l��z�9�O`�a�Q�#�]��t�f�k��Q���CAf�8xeg=�ij��$j��$��AP���>����:�_�Y�q���'c!�5����A.��h{����*�m��5�%qf��i���~������3�?>����:�ؽ�2�ϔ���B>i.BF��;y��������2yM+n2�Bl�g6�u�o��rd��$���
Tx&<���A�>FäL]j��aJ,^��n�W�FSq��a��lgW�w4�q�[�u���3�������aE"{3Y������������+N/bQ����ܴNk�Z@��D1�quc �3�xP��Lm�����/�_�
���8�jHţ3����8
��ux�Uz�R�aa�*��"DVCY\G�����B��6L.�F	����9v��S�}�mj���0?����W|{���d�
R��<�0�0k��#8�N��x�i`�<#3}P%ENO�B��{�(Dk�/)����7X��Uei�DR}��� �W�xޓT���D�;��x~_������&��<:��ʭ�N"�4�n�f�AГL�ڠ���]kЪf��-�m9N�-�k�.��3N�g%%�V����m�혋f�2�̹��׿ ��R���glǍ>��V�	ˇ�Ѥ�^>md�ƶi���o/����3Ly�B���Z���l��|a�J�0g�i�`L��J�!܁.�G�f�Y��5���>P;E�b���r�����<�o�o)�#}gb�hŹ�!����1�(�#yk���O!�A2[�^��W�)��ҽK���l��Jc�h~�`��e�4�R�:���������ՇP��/K���A�#<��h��SZ���ց>R:�kaiC�����*��_ڧ��Ir��;5����)��t�q5����b���_��fM+��~E�:h`��4�g.�lO'!���242/I�D�������{I-|PӸc���#�'�p��T~��Ď��m��菴����T(@�.R�"��T ��C�kg'7"4g�Y*d���ؖ�#�w١��<�PÍn�̢v��~C�N��F����t&"#��D��խ�,���$/yS�O�y��������>������;qp�K��(Bf_���R"��}AS��i�Vr�� ���!���x=�u�����84 �����O��� ��u性&��l/�-�ʖǉ��������`zr㫩Rw���F��'>5/]�;�N[�~A���T����j�G�s(��Rp�H���&��2M&MQ_�[΁�-���Z���Mf�:���dN:&�]���~E��~��m�������d��Z&[<��$�������,l�9n�%��AXƒ�f�A�'�RV��,��9(��f���z�d�tZ]��Wp�H�y�>~Ml�ؒADjw'Ǡ��`U>�i�Zb\k:V(����BXR��{�_��6��1��7��I�>�~'^�^X,���	�,ej Y?]�!�$9�4.8���tٷ�yoI���_�2��#iDr��\N��o�N~���P�</�x������[�؞�!,�P3x��u�M��eG�۩���e�9j��%�bwŻ��J���@���H\W��=�݂�>�D�>�D4%�ѻqo�J��&��6��Hg����0Қ�.���w�\���:���(��e�ڦpU�_`�R�q~�
�r������������[�3{6�)�=�4h5��*��D$F���j]� 0ȣd��HI�)pB����)��n|\�UX�c���7s�EC�G��ʙ�)Z���9��'dgLt�|�`Е�_�T~R0=?y����B��n#�'�%���NW���Rj����U����Z�ʁ����ğЯp�@P5��D�
D�1�B�$�����K�5�7�����2���+IU8�F�N��^��f�Q	�T�hd���u3UGk"�ª���`2��==75��%7(�]ժ�['��n��l�ؾ����q�j���6�ܧ�l{ݓ#~�ͫ����t�\�A*}��1��8��U4�5�
�tFG��C�@�v'�Q�-��d�vKQU��PC^\J�^�y]�	`D@�,�´ �%dƿlx�,��h��?Z���n��i~��L��I�?�`��d��EN��l5��689/[G�����Z5u/|��뫓F��NA,7l]�r���~��n$����g�	�S�OB~���z	��?X�����J}<���ğkI$�Ә�<-�����hM�- �f�0���|��~�-���rq �,���;WK>���|L�1Ah�CT���9�?���g��Wm�v�1"��Z����W].sPu'�~C{��so�j$2/�;����,��4wo���D6o� �]��&ӳ��a؁&����2���6 �r���0�����E0�����j�h��U9�[�	�k�W>֛����DH4A�/��G��[��=QW���u�.)b�z@Z���Ի�*uD�
tݱE��3o�G�h&��T���vI��'��)3�8���o���J�	&/UU*%��뢃��O$ݥ�uNI���<$�S�t���2q4��˥~����Y��0�yB��?�9<l��[{1�{#�V	��M���gp%��",�Sh��XƎ�O����O��y}�9r�ҙ�q��̑���%$�q=���#�~������V$(x��KS�Ee���X���@��/�~B6�.{�\x�}ip#�s��I֖���e'�$V���z�[�q�̰󮍇ѿ���D��臘A�����U�������b��B�.l|<7s�"�`�%� Gk��"JF���:5E�T���}���=E?�kPoq�<0��K�%\6�Q���3�//
��GZpY��D������.h��j�j�œ��1����dy cƚ��d�p�"Q�܆�[q����P�/�Qp4&��1�};�D#������Uw�bL.�Λ�b�`ES�~6�(����b���L�9�g�����&;|�r�;�������M!�-W=
s�u �T�*EE.X���ǆC��� �(M�S	~`�`;��^� D{����Ђ>���N�ز��fPQ�pn��xx�~&�_��R��l�F�^x �ΕW`�<{���,���['r̞��Ր��)���d9<��m7���9uד��1e�]��� �g{�\��W��5+�����7!�0�nmS�u$)h�֘#p]ƑR���d����<x��{�X��5��k�`���RP�I�����X;��#t��z�T3!EZ���ذ�
Q�+P������2�4l�gn��%!�l��j��@��U���{k��j��1���V}"œ�Q� �]��,RUR��m��C� c(�f�9��&�,�������F��>8��r���O 2m3C�Һ���4	���码�ι/��y����m�C���N�<�s�^�!�L��C��W��5+���ĉP�i�{�}�6B��u�����r���������G���#x�D����}6�p��QEy��T��t�������D�@pp˱��rR ��������2
�â��Ն�������L\Tb��L�"D�9��w߷����C�nd���UB��]0஬{Hs������h0ٌ��5�KO�d�D9�M��^O��;��=�{�׶��d���++��H�z�/� Ҁ�D��B��-aƼ}�5�Юf��V*ܝ$��l��
�{�Bk�ߌӉo� �û"9�Q�I�Z]YX��{"euG2��ig�3��fI���|����]���gO�M�8<��A��������ؔ^M��i�" 0E�YJ�_G�t{4�N�vK��?4�v뀉�kE�!z �����ۅl��GV�D�b>�GF6v��j��m��)k�����W	��K@�`��Obx�����2⸴Knj�Y����zA��cA���s��%�����͢83�����&_h���zE����������Un)V�����]�ܠ�
���E�0���-�uy�VQ�QVY�D��V�Ԃ���+���Mf�L&��	��9P��
@��+�OF#�Lfor��&> >W����qZ��:�L�_u���ⰱ1$a�1��J����&���5}S[�o2�Q����G0~|�9�$�1�T�:�>N�`;2*�9E��N�A.۽�D���v/�p��.E+=���{ilݕ�W�#����v)t���rIUM�p֦��#:ʱw������Pg�rn�n��V��>��0ځ?��5/���{�^��c�W�F��$�m<�ͨ���Ku�+�!����Р��އ�@��KX5����#�?�:F�g�>��H�g$T�h�hh6{�]ֆP���6��P*7�[��M�cƀ�L���AU�B�?��WL��U;�O��zڷ��LG���
}+IS�ݛʐǜq�Jm��:q�o�H�!8�Ci�n).G嶾�K��DDOm*�W��W�S���\��_ALw��S�z+�[ZO:0B�YW�ޝ�� �*��48K�s�	F8Նv���y�����iL84�T���!P|��X�Wo�뺐���	�{�8���/�;��T�Q �Sr&�`�B���&��n��ΰ#VV؀�o�ȘS^�]� ����yҕ�.@sld� �ü��b"i�QM_6UA.�����1�Ф%T�<DS`3`���_F�g��-��)i)�ܪEn�I2��C�:D�b�N/ٮ�6�I7�ˡ��%[��Zn�����*u%T=�&.C3$=!!���7)\2��l��Fb�D�}�������m�s��+	�Z��-�¥�Mws�U��X�;���k��ؐ��Ş7�/cҋ��vAѷ �>�� s�[�	�&P[p�&͙�:3.[����������d���(��!�{#�W��U=޷���Ҽ������S	R�u|H�i�4�۵�)�����w�}���^�Ϩ����0A����y��X��G�bKZ���W� ����r޲ S#�j�r�����â?��=g;zP��\8�>�:��b'���4���U6s�]G}y�\�4f\n�:I�kb�z:?�s��ț�f^�����x�����;�ڽ���Ne�YA�o��^|��76�����E�"�nWڵ^�{�Z\4׊�@�,��I���ޚR�� ��:���4��o������3�M�X^��
��t���)����M�3�Rw�f�bD�A�������lC'V�Y�����*) �'�ɞ45*��E�����5>��E��ʣ8x"Ҥ��S�����%O�Aj\P�W�st@� �.�A�;�M��G?؄͉���sW��@j�5͉n��n'�<�L�gg����uCa�X)&��,���[*5Fn?CR��E����4+%?(3W�1�-�m΂b��|zlh͵]� �<l��3+t�q@7v���^��+���&��s�/�d�W�ҏ��D�I�<��Y��Ɍ�ծ��M&�M��P����y�u����e���͉@-v;�`�����O=���ǲ��.�8������N��q��A7mְ(T�w��ލ���8uH���T�]�e9�(Y�"*����x�,=�ѵ2��dW�m��@��Ho��
܉���.���oy�����3D��9�M^�*��D����]	��� ]��$�	�
��n��a6�3m��
�Ţ����� 3�F� I�Wu�R�ȥ���p#G����Oy���/�#R�/��`oYg��xeL�	��D��=���P�jRVK�h�JƇS�'���gg��:�؆;��A�x����U����/�c��:��HX�=0��i]�4��~�K���y�h��ډ>%��p�Ԧ�6���s�?w�)o#�*�|�_��}0�m>p^bR\N�PP�={{U��IQg�^�/�5���Q]�՗A��RwY���A�<�D�Ŀ���N��;2T�
*�Qf��D��I�7�|\4�(��+��J颌�2����mB|�H1���}�I\���Ms��1�ⲴEfxD�*��?� ����Hm���]w5^
�� u�ׅH�,���N1��!�	I��|���h�7윘I$�P������:�/
����p 
e$Sx�	s�|�z@�42(@f�K�>���i�8�aJ_�c��G܍n0*!��#���f��-Nf_lefw���kn+��߸Z�H�8���|����� ohm؞��?��C��s-���d�7�칈2�BJ�)�hqO����E�r"��C�!g�9(�nډ_rѴ�i��<D�R(䝪����[�	p�������!Gt$(�z4��qbJ�>qA�ot9�G��Q������ƃ6Y�9��67�6e���@q�í]*�l&2,+�ܣy��j,UA<��Y�J�?�Vx��f��@�����[7@n��"�&�2��3* �i�����Ш�EE�bwh(�b�-���ȝu��}L�$��VSD]Ez�R�,��!I���
I/� 3U�ad`�|�ޫ>Ⱥx���J���&hcA��;��r1���N��D��ޯ�"dM�7���1�[<���w�r�����S��ۼ`v�� ����/�4jMa��Z�kYT��T/]Ӻ-M'g��)C�f���!��@
	60�y�9��i����M��)�J����̶�rQ���G
Y2����q���܅*"qF��w��1���m�`k��D��8�
Xq��Y�t�����<���=Ƹ�w���$�*�Y` �}����n7�h����<�k�0�.!'/�翲II�p��Bx��ۿ�w�DIG����sA􅠞*n
�ȩM��'DLA�R�ӥ�1󵕍�u����.����V�Z�+)�9
���y�9.\^ҶM���f�F!J�V:+�Д)���SV��Ɇ����^X�FԢ��c\GKQ Y���������&�vD�'3x%�9��ϣ��q��7l�:�[Q>x攑5D����·���V���v��G���\V��ǲ;��4*	N��~b>�#E�Q�	�Ao�1m���A;ż�Ft��0!g)�N�������қ�w�N��3��>n70l��e�M�u�&i�����0i�!r�L�C�ٿO5����g�<$�S�fgU��k���@��*�@�?�����n�S
!��_�:/0���"}���S0�'5�>rr�ec�PhET��̱��%1���Bq	H�-�m�}rA��p��1���RNjV�сJo�`�7�(�C��j�`��Z�#E�Xu"�ŝ��䡦?�W���`���	��aqgʉ+n	��݆E=-�5j�K�>m 5<>~�8SH���̯yq&9���.�vc=�bk��ESc"�[v��8�/�mZ�#�8e[4@�U�q�w�4��C������Σ�l^G��A$���J��	k%I!��<�^��>����%@� 2�k�Ň8�Y^#/$wu�l�����AJe
Jo+��T�W���0�G��&o�����i�ӳߋ��Pr���pl�zG:��@Vl�nИl�#�l���#�zB2wF���Fq�HpBOA�aQ}���ѻ,�d��Y:e�:v��~�0zOm]�R��2�����Uy����{�M��\
��;�E\�>1(�ec�!���+	v�n����Q05��w�Cߪ��w�k8~G�S���v���p���5�/'L�Jc�]9��K�bo����0���>d���M�ٳ$�0p�1��)-�����x��n���3�q3W�\B��R���k)F���5Oc
4Hz��A��1z�w��^��)C�:�� >:�:�n�Ҿ��wF,�s�~n�妗nhO�{[C�;�;��r�jJ3��Op�o�=�H��{0z�FS�R�B0�kn�n�_��z�1���ڴ�r�S>��Q�35�#��#�n�&g/tH�aU���������rgw�&��&o~PK���G�)h@_n�������Y���N���u��Yq�}>vQ�M�ŶI@�u �^�B����w��*������$~�ݿ�)fw�	�?�����ފ�4%=�Ƚg��%-y�
>�ul=�2n������җG	��������:��3%����L�.���,��,���A/�Z&�F�>���p�Ґ���:Y���G�YX��k9�#�'�fT�(|;TT��>�J��E���y�/,*�╍;M&��t@�#^�vH�˳�՘Mp�%�p��UvF��憋�U����+^Ad����+��(P���-����4:���zB���z��
�?����("��Z;�O{Ox�N�r5���-#[�ey�%O�
q��vî�����gwn�M��*a�Dߠ0N���0�	2~/q!r�����r�#�����L'V51��k� 3��Į����Z�%l�mo=�0����������Cv�q���.���"�ESޝ�k�����lgG%����ry������O5� ��F�9G���E!䘇�96K���+^�eX#2+�����a,uFt���;�y���}-H�֩L�^�B�C>�ْ��xB
�����@�E��[S�h7n*�S�<�@���8ș�X}ٸ=����Kz���D6�͙(d�\�e-u���.Q��U�3�jnk��0�s<��ϛ�:qu������w�'�v"����#O(�z�y����\U�B���� +kG���Ru;�2ƖI����ƏȀ-�(˂��@w��n�[ 6�ۿ��9�k���?�E���	����R��l��
.�>'<�L�2���������IZ7qƐ�/�~$*M!��: X�S�ѩtQ�TR��}�={8�3�w Pv����Qm	�������kx�E�9����o�Z8 WCml/
�`NG�������\��@�:��*��(>��M��8�B�Cz�/���s�Z��D�����W��ǥ���-z��%}V�(�s|\��[K>jsiG�H�c8���Db��r�&d���1yD��*g��V�ӎe5����YèRd7E9���Q�_�F�6�v��MFl=j4>�I��<���8^�im���^5}�Ӥ�ɑ쨘���f��B���D��&�ŉ�o���\<gW�۝���	H�pd�HV`�������_�B9��6ʉG�|~��L�&��b��#,{F_�V�'먂�q6��L3b*�3�6��	�T}e�C~z<i��rw�(7(������?���-�7�[{z�b?���B�t����hV�H�\Ƭ��F������kZ�}�0�TUϵlF(��ӭ�:�$��n��^o*��%�*��G�#Kq�r{��ުx#1�I�UIN]�+xϼ[Ʀx�a?�Z�I��2Ў�'�a� ��n@�����j���7Y�p�#Ɉ�C����ʃK�����]
�v��eި�Ͳ}T���}�ng�VI����"�����(�����Bzd�+�A�ӯr��,c����'Ͼ�����X�缳x��LU�U�1E�����k"D?�u�I�fAǦ�"ÿ:R6@�+P�aq<h�Y���C�I���	�ΙG�g�_6�ng�˿����X�17��&Q	^�&`����40�$��Xv��ɬ!Q6B�+d���u/�(�Mm�¦g��l����-�-���:���$��bE�ѷ��>/-~��8��ȧ��r��Vv��E�^]�]L�bȈY7F;�Cm������I��v�]gv�HD>ﳵp�Nz���ܣ�4}	Y9��~_�=FL����67C��jGt�T%`P'��Į�*�a)��p�DZYK�����?zO!C����'��WT�-I�$Lr5}Bb����0�~Hyx� w]K].��e��)R�=j�ҍ��D�(�������;=��7���P3u	먝:2#����h>���v��'��tx�m �T��ԅ���w���A���m������|��,F Gm�m�t��q��%�b��xb̵����l�S���f�3曐��{M`py�p���0�_AW�<銥�f�40����Nem�än9����0�<;��������go��Q�oH���MT���ˑbK���:Ћz��xe�R�bح�*>pAY=Ĺ}u�x"I{��P��`q�գ͕��fQ�!A{�Q �0CPE�,ϠX�Z�qX���@C_	�TqR������8�VW)��:����=���}8W�O|�
�Qxh��%����%��i��aO�����Se��3ab�?gP!�����j���`�	x�G4�1	G��QT,W�Y̑9� �&��?�A��uw�6��S�>t�bT���H0�0���v��}��7"�N���d��gP�����������8���Y��6ˌe	���ь:�Թ&]+��ֽ�o�+==۷'�7�~��g�'�8���d�j��#눿ME��N�9[>-2��A�X- �YrBZ![8��Mu4	vJ)��&�h9��up:��Ṟ��r�5�pc�d��G��S�G�Z�����gP%K$��NV}�64��[)�NR�=�%��ʐ�"��f��v8%���-/�1Mh��ӭiB)�H���l�Ԣ����_Ř8Fk=6;��d��|j
����BV�f���\�li �wXn��2P�p5��"�\���T��$LH\]W���qV4rO�Ss�{��֋k�u��AzG��c�W�'�"�Y:�����~��v���:�AX?���d�u�´���,VH�X��� )a .y*%{��n��t�3w_���Ԫ\N��I��m"e�b^�Ϸ�%��(:p�1Jb�g��O�����T��7-�0	{�%��(/a�"�g&�������-���c�Qe����-�hB�����>PFv�'
�����8�O�xB'�K��<x�¬��Շp
�����}&fy��8����fli,(fn��7F�������O���h|2Uv�iF&�v��9B����4]�������<�w��C"V��%�kÖvL>Ą$�(b�]_�[��쏫A��+kU׶9^� f�&���������L���#�5�p�����T�e�k"��p���K���#0c_��6�h��=Z��.�6��x�4偐��eE��b8�،Ӏ+���eH9�>X��-���V8�j[kK:��>	���ZP5>�2�U�D�.R������p���~X�D$i�`1hn������(�g3�t�iΠ[$����"D���Oė�	��=4"�]b�X&Zܿ��V"n�ȧ�*�ݲ,]���B��,��R��E+Gwճ_�n���q�3�is@s�њ��� �j�9SkU���m��q��(e��]t�&.�R5��U� ��λ7�C�L��M�y\?h��L��ł���}P��h^���E�ؕ��P�8��襂w�������D>d@�meT۱�ٴ�v�f�\��`�<T��;��/�)���4���d{�
�D�?#�[?����5p��%��*�n.&k�3y����-��eJ�]+ >U�[�w���^=kQf
�Z92�8w��X�	2Dx�~c^"����s�&�-\!�r�^� ��<`3��B
��V������;�I�����J%��xc��b��rv2�c�/�}�&�<�~�G��E���n� �S>��"����k�7񼂚U�
Q��<XP]PD��4�ߘ=K�(�Պl1�_Y^�t�4U��/�<\x=�R��A�<��3}:� nx�3�єq0NM>������`��#C����� A�@?6�zk��x[�(�U|�~�����))���sۢ��rRU}�iq7PcsD*׻�� Bqb[����u�7 �$}��h���g�<��_��zuc��HC�q�����6;�0�$?&)��{܏��,�M���a�����wEG̵�xiR�ղ˵
�껭v���x���[:�IG���ZZ0�d�t�jG4n�Y�ʉ97_����!s�E��it�&�TN�Đ鎞3��;�3y���ʼ�����iG��;>l�%���?lZ'�|�/�bM�k��I�%���tCB<��qAMo��Ԕ��:M����&�(A�<���J��/� �%y�1��W�m|D���M�g��)�q���ԧ{�1���([��6�S�MyB����ޤ����޴u���Rr��utj���Hʿ�%���^7�q@��5u����q��h�I1�ZG�聢�}Q^���߸�Q.<݂a�`��2��5��I�Y�_:��$�8&��.��u���6o'䔇Y�$w���������$������J�z�=�&�m`�N:&�kB0�����˪��?�4vQ᥊�[h@��������氚k^�ך��/�a��]s	�DY�>fd󆓵ز2�LW���pH�>�?�����5��5K�V�?�Jܰ���$2l'�ǣ8��!�ۣu���=W	�����zp�-'^d	����iiB����:��~i�ٴ��cޡ7�[���ηlo!AH�}%�a@t�U�a�c��K� *��1Y[�����S��j*̍�^v�[w�~zMg4fqT����(�f��PG�����"�Q���T��x'$�3����"�q��8JB�"�b^��s�)�y5n��ｲ�zIK �lΕ��wJu�����+p��Ɓ:����V(�ǄbD�:�hy��A��6� ����g�QV�%'�o	 ��Ac	���S�NN��b��0����5NR�JH���u�ȿ�tH|�U;��>���^�T��&�*����6ݨ���"Q�Ŏ�C��/��'�p�z�Ԡl+�Y:��G �wd\wr��OF$ǥvG���1A׻B�+ӄp�*�3wA��]bṢe���d	F�`#2@;V�_t�on�z��R���'���.�v8�N��V��\�h�m'�	+�[S�Q������Ƅ-ys&�߾Ia=Y>C��./?`� 6���APg1�eP�FIw+���sՈ��O��VD�t׆�蹵I��1��Hu��!a�L{IFYK̲�G����+��_���2�B�?�[�,fa�D!B�`��4L`g��IPZ� ��>n�j��i��6(�-����i��m��X��?���M��x`��ҹn&6.���l+�@���oGÍG}�����3�<f�����'��
��a�X)M�㳣�*<��ēlj39W^O�_N�B�z�Q�K��8"���{�O{Yk$���6�ȕ~l������x���D?�������!�$�k�I�Ö��I��둒�x
���Qbo�������,��&�j�*b3�5)0�Dd��Z:.<�M&P008��Y�M�۳����ô����<?�z�
�E�ͳP�lur�~�J��αŶ�S��Q�)�Z a�H^��ic'Lk�a��!��JB������3�yh3~��y�K�N/�����An(0m��$��)�]�E3�x��_�*`|aDV,b���m?E5�<풵#�>
�X�i8��d��WHzZ�~��ŒeӸ��T��Ԃ��Ԉ�d� �/�4Bq_�N��8�/���QI�15�)i��{��˫�I9	:Of������'�[��.�!����q+~�.�be�[,1Y����cJ)X3���Γ��.x�"m�ɮ��m�ԂX���N�X�R��k+I>�F�m{�.�v����b�C��A�4'�K$l���hm2�(���}%L�O���ณ����=d��W�j��B�Gt�"K��?a��R�ڑ>�i����"���g�!-� �شލ�1
�\A�a�(�����������L����>_(�>��<|_gt��K����l(F-����~�KZ����7��`=����x��Y�-�y���~�x�|���_���S"e®�^�ާ�%,��x���%�TV$��Yή�۶,2`��=U�8�)�����H��2ħS���l@���yw����dV�	����G��]�#�+;�O�P�Ж�����te�a��?�8��|���86���>��j�v���RG�W���\ڎ�@��ݮJ���I�d�
Z�s���ܵ��K6���s�O�ĕ �O#�l�X����wH^���-*�:�K��؅�)9�O���������̖p��͚���+�����G3�i�Z�F��zcq���p/�`����c�����X0 4l܊+C���3�u�2N�=����tL��P.�c^��0B��M��8e�<˱H��<bO/!h����X�z֫��X|��^خ&)���U)5r��)Q�+��=�6��ږ}�N�t�m7�?��hW�X�i�A+RF�gh���M �w?Н�c�9	���(����um�0/��(4&�R[}������.	��x����E��"�cƁ�����duO�c�{�Zi[{���P�,ɪ�����ц����$�P�FU���Q����9�N(�$��C)"�q9�F5b	ƽ���N���KJ[���Yn?�@��(�H ���Ϟ�?���=�|r.m�����'�Gtb���l�|�6Y�.>�1������\�5F�;$�ٜ�;�x�Bjٻ��>5:�����|Sl��F&�̦�s��@�ê�f����q*�9B�	z�D��tp~bt6ur�&!��5���<��p��-6Q��SŶ�k���<�U�Ȕ\�ggƠw��黼����z�\1S�ʌd��=��5�f�/ǒ>d'Ek�C���d�h��]����!u*F�q�)]Ϝ˺-s��?SHt�]ė�t�Rρ�_�c�h���C�{�t~�z��A��@ί�}�𣧔�#�����}2�z�����c����jdT5�Qɏ4U�ҞS����ֽ�E$�5i�o>�1��'#c,�ێ�j&�>Ot������ɰ��=ZV�e�5� ����Gh�a�Tx0�qT/P���b�k`���z�<�'�#z�>��Hamk'{@rSP�0��m�DiK�YF�s3��cM��Z�)�����Y@�m����rB]]gG��zv�&Q3~�b(�Mi��E�X;����}CJ�~U���P��7[ڎ���؆4C���a��K�����|E��nWV�]�l�#���1�4�:�t0��^�t�W�S҃�������_�K����w�_�֫�����vئz�7<�/�`��IT1R&����FdQ�#���L��08X��r������`�8��b���J�w5���`bP
��Hw�fY+֤ɷ�s���t����~[c��K_$�x�h�Ҥ����<$�\09�Q5�$�[�~2��8u�ї�K��;�U���d�T���I3��������x.��Ao;�QF]=|+�&J�#H6���1	jSk���j[be���_ά����κ�?SY�
j^%[�_ќ�Z}=}���	�,j)M�YiTĹ��3 ��i �0���2�n!#t����"g�}��hC3��@��2K���+�kࠫ��f�U�7>�K�����_R�o�$罘�(C�x*?8C��ߞ��Tii�Q.J��w��3�?a�FޙR��E��L&���zx��},��:�0ʉ��E��W9\/�n6�L�|��J���)E
�,G\Ε8�nJ�c�g��?��H,���7�����`$��D�<�(�s�t+j{n���_b7�l^A�П_�y��0�e�@���w�ItW�oT1�Heg����j�y��T�Ѣ�����@5��Y�1�InN� x������l��-=��V�F3�d,� �@sf�8�{9�2m�L&H*_N������U��vv��V�m�D!c:͏��#����+L�C�%��
~#�S/.�~�"�987���6su��n���S7�b�a�2#פI��:sXێnU�$�9��]}1J�ߦoQ@�[���,�����vA���RNxE�s	��`W聲d
�Q�V��/-��U�$��y�+�:A���l�tde_����7>�2U:�qy���ݓ�=/([���E~�c.��j�-�cZ��o�rS�������?�F��jG��b���U+{����
D�"~D%�<����X�2��Mq��KB@�u�e���l*�ǟ.k����㥮O�N?� �{-E�f�@��꿍rn�J�К�p�S�u'�:Q-: &�6��+%��
Z�]H>���UH��(g�-�Ye�w��T!'�/K�r���_�	'W�0�_xǍ ���]�xR��	��4���f��|"��Z7e>����
�d�~܋U�qO%}:��j1߽��z�ڠ��	c4MMeI�[6�f(ۗ��f�ZAI��O(�\�}�T��k���;0^b�O�ZLC�QD"�&��6�$y� 玆����{�e�j��L����F�x�K�/�%�!k��2�YP����L�wq�[i�I0n�r���72�8��D��k�+A޿:����T>u�c?�5Lƈ��������O� %b'h�j�Gnn�ߑ�.�
RiP��j�;Q��~qM�Sˋ�k{���N_!���L8�zI[��}00j�R �?K����2��	�l�x�l+��0L2a���d��Ǽ��$�� ��G�g��\��L;}#Ԣ��E��C V���<p�����ާ����Ɩ�~ϫDm�5պ�y��Y�h����e��U�<�6�P{0r���c�1J]S�A-���PK�Ji\̈́��xU 㷧::uϮl��x(?S�R��Za��6'�n~�����W�i~���n:��`�r���C�&o�r�4d�l���-�����N��^;�mp�Cl�;�e�x������_>nNs�P�DV�]<�>�?��.]+����M�G	e[�Vٱ(Q$�-ҦS�z�mU�jl'��xӌ�>���K�N�uzC��`�M`S�8�rܻ�zo���t��~�ڪ;�م�����t��R�;<Uz�hșӊC6[�vT�#l�]��H;����>�1���z��<�*�����6/��S��8����6�s��� �946�+�*k�RI~�Y����bD�o<�@{���3�9���6g�Z$֠�F�)��ܠ��N�F9e9H�!Ѿv��%��o\�u�$���:�����ɲ�=������
�qj�ϸ�d�����Qn�{��<"���19�/�u�lT�.\G�"	T��v�T���
9@�r�X}�'��lJ���9�t!y]���� tY�t�L��f���rs��ݨ��sDr!�E�]�M�������@p���JZ^���)]m<�]=읺K�g�>}�����P�p��.�Ǔ�ތe�w���1!�w�x&m*Ҽ��^��襯+4B�?N� k�P���i�Q�ň)��/=A�W��]���5p�놶�(��mb��?�D��ӆ[v<Dg���%�?R{>$��5��=SXV�����r�>�VGԘ���8%aj�y��%|b��U�}T�p����T�ی�$���֦��j�x�
��;�.E��<F#�pJ"��� O�2�s$,9�¨<���D���\�:~������p����C�Uys=v7A��e������5�n��$+�m���g��Ų�����a���h������xV(��YI@z���uGqp����"������Zq�I�$��� #J�:´�2�!����_vZ
��*+�����T45$G|��V�4h&�rb�����u����f Iڻ���0�wf|cz���
_8�RdSӖ�]����uSH�]�P�1-+�g�G�Qf4M�����$�Hvވ��Z��G����U��<3+�{���K
<�R�lo�)H�T�M��!����O�uHy��I��j?C�I���;TT�lΌ�ť|��yڿ�Et�q|EY��,H�S�7���ZNG�0��7tj��WU���*q��Q�iK@�l��UĲC����W�/�H+f�R���C�ǣ������̅�p,b�� )(�M��[�ɍѐ�� �W��F\f�8	�Z��^��G�ξ���u=���\.�]�{6��RocېCn��D��5�2�H�� �J��V�f��:�����sB�,�a��S�a��#e�d�����_-��y��@�,?�t�gZ�v	��q@�3U���6oi%#|��ɍ$��{�΁��`����$��Vq�(�`���J���0Ҿ�;/cW7*{����u�+P�j�}u2v�j��M��f{���+k*��k�N�l���0���s:��ȧJ|��uh�.�l1\� 
fB�ǒ��ן��Bo�zI��I��dS8nt:!P;���ԗ�����?k�QXA�D���K�H,<�����ͼ�,�m�|@�L�]ڞ�>���8| �.�%�
��K�;��4�_�N��GT� (إ��4�s9�!
�A�k?BfP�ܵ�v�C��R�L1,�%�ow(m��~�u�����Da�t��z���{)��B�<�	�n���$� z��T�ҿ���%
(j��Q4���亵*r�� ������j�D.�h��J�-x[��J(���p�γ!�r@�ګ�]�*ʨ~/�,����1ihU��jQ���r���	�Ĭ�EQ��0�ؘ�̯�C��C����e\��rӦ���|��<�/Þ���m�u��Ա�
�����Yc�k�ܳ~�Z#�w���$��T�r���$yP9v⹡�?ⲿw_��a�@��#p��.����o����H-�jT01�(�C�lE����Vw�9�tgJf�F@���siB��O&�΍+��1�����"h^&�)�jG�H9��B���?����(񰟆�L�V��k�R'�\������R-E�	Ð�-��k 0-kKU�b�����7>��ԎC�o��=�ܲK:��`k��?�I�����F�k
����;��'�̾{5�������0�$� �F���Qǚ��[}�sg��R�g�� $m��|^�cXk�tK�� Y㮤e�"�[S�3Jr�){zr©R��`�F����+��h�YX��C�5+��/?�$R�2	�������}+�`�6�����Kq��(��H7���y�Tn{'�S+ah/Hl�J��F��n�=��O�O�[�D,��ǅ�G�5/��1R��^�ǅ�be R�B"U$IHɠf�p�߸�>Wm��ic&�f����y�ϞC^�x�S�U0�|���	G�d,B��x.����a�|�h<�1k�ՕZ��v_g/��Z�~@��FD!�8�,*<�-[ {�R�щ��9����\�i�b�:�w��HU(��Y�ZnO�����c�0���t;J������b����zՁ��Ց���m�*���F���O-m̓Pڻ��P���~�AQzZO�1����@�X[W�i)��h[&�Pk��|����N7wu�}��p3��͗$-�k}���|�w��E[�BǪ��uI�q|�!x��D$g�e"�5�&nNQԈX7�򑤨�I��8�D6�v0 p+M@�B�^��.�4�*���z�L��L�.��{�퍰��;�i��{�<Z�G��ki00���B�e쉬��A�_����"�:- ����w`�v�7A��v_���q�(9*�r�f��lg��׳rJ�^�����	��E+FJj�Qġe�q�_�����jiQ�h����lj4`O��B�~��i뽩`�$�d�X��B�����D:�/�E���g�`(���K�&--���֗�}���x"��W�/w47��ac�ե{��4��Ej��������_D���`����Gl�j�V��|SA�Y������L�`��҆c�����bk+}^B�m����k�V�g���Y���$��~/�V�T���Y�.�>ߗ&MV4x���	._�q;�VG�~Pw)��@����'��A���J�o� Վ_;�U��Mg��M˥z�qv�h�%}W5��H�|���כ�|H�q�#�Q	�m�-��̲�3<��c֙%�����fV��O�ذ����8ua�8������]OsPc7Ǒ2�BpL��u?��;b���G����i �9����?����:zRUN4�OYC��7�'ZI�vk�5}��+/�=: ��A�y���͊���s%�	$����rS�Vn>�����E�M���_�Ś���G�T��l� Oa�����s�{Й˼�7��#�6�.�TLI�?ů�(���e����2�v\T��'�g���!C��</�dyŠݣ>���sA�،�&�x:q��:�L���H7��.U��f2�����l$��K�}с��8�'ϵu6�������9�M��wٖ��GԶM�y���aOM���'�O�Go��(_��X�1�)����'0د�9c�:��S�D�2�B�-&�Ρx��/� ^<Ϯ��[hC*p��<�D�w�b�L�l+d�P��U�&��W����v�����.i�kpw+⷗=�&�
0�U���D���QA��0F�۲q�I�� �.p��<�8�!z�G
6L���HBr�����g�a$]yޘ�׍����$��o�棉}�Xn
���aT�8���~ۇe���|\C=39M���Z�0&bd2�cW�_7ǟ'۴'�g߬�Ѐf��XH/�s�?2��&�0�f���DA�W떺?�\�������/��۪"�� ���}(�˨ޮ�YO�D!b%��?'��G��q��B�!��b��4�ǡ�$�=�Z�3�!�%ʇ�Cg`���U�u�Z������S���i��6�5�1������W6߄�i�'�W���<�c�[�%j97V�5�ڍ��n�^.et�5��q��ݼ�����h�.�?wV��F�=�2��|��ddu�9Ps(p�ҐC��d�y�K]�#���~nn��(4`��,YS�zi�t��QjD���Z�.�/}�v���" ��ܼIs�Z�E����7ݹɘa��g.��	�;�tS�(�Zx��k�Dw?[�����e�q�{�gg@��q4���<uE
o�����l���]���B�[Y^�T%4X :'��n���/]�����x��N��Z�㿦o��btk�{'�4�������Ѩ�tC�Lܾ%��lt~�p@/ҧb��&��t�̣'Nn$����W����F3�*0��gz��U
دQ\�n�,���%�a��>v��	���|�O}�}���{���I�=�?-ё��zs���,���c�x��$��w(���iVͅH~a�Ur�@w�T���� ��+|]���-����E7��&%�]���-%���EZd�����=�L�i��4�P�2H�`���7��/h-4`�P<N��N�@�l�吏k;b����˓Va�	��������2�|�υi�јHI4:��/��c����	W�� �U�k���3{�����X�õF�x�_�{�����j[�f��Դ�������4X�M����F�Z�/0������z\��FF���'Ň���4S	m�6U
uj�o�TN��v���F�����O)����KF����ׅ�:P�0�ٍG��SLĨ�f���B�wu认�:�b��(F�]Ij�� ���ۊ`�s6xrz�b'�r��&懠<wa��i��vv:�]�o[2���� L�!�
"�à��c(����o>.�`&�l������M!�&R���0��qBx9>%TX2���Hy�z��r�����ܯ ��)^+�ָzfH	�"��F���
�V0���b�K<��V�=�ʬ��{�ٙ^w J1��d�"�K�?�!;�}��VX��Y=/��m����/�ÑZ���@�t��?)]ؗ�����"������gez6���}f�|H�k���s2Eis�N t��~��[i^D\ �0"�|+AO ��̬���L�P#��L�6 KH�ض{���ܧ��R�1���?-��a�`�>b@+.+h=E�m�##{�!=�,V<��"�V��ۮ��n�&Ci���嚡��?G���!V�Fb�2b�M��.�S
o6�F�dk�ML�(1�������{�'!b�l A��X�]x��&�=�� πv?m�c�lTa���}�5),���`e�1�6HJ��f',��Y��4��}��2n�D��k@HY�a\�G�C� �{�#U\��@��0���a*[?�i��zhؑ[ �����4H�N����̺9t����O`#Yl�	ޕ�P�	%=�]���0��FxԠ�4AI�U(FN���c�7c�`6�Y�$2G���|�ƍT݉��6vh�z�x:�`%fV�x^��T�^*oHy��,U�t�^
�WgW I���6D #�dDf�X,���&�rD�ſ�j�O�P3�"ʳ�l��c\w9+��j�4��ٚ��5��q�_ �W6�2b��da
�����H1�״ v�w���6ظS���q�H��;XN�Ʋ��UcN_�:���x!	�Z�#Y�+y���&U�a|��[E񃑽g��C��wY-�3G4-~�#��b��5�]�Th�9'4�ߛ��n'�Aa�o��������Ԗ�?(gD��V��\�vs�i#�"�<T�D��b�K���d͸��
&ܟ�c}�x�
�!�*��X���v����;W�Z�%�Rkშȥ�c{�MȂ���^$Ue���������T��#��n����J��(0f,��<]=�@/�Jt08lB T+ई���!��'�%npX.��VA�[�:iu�LI���>u�=�IQ��=z�*�������]�/��]������d�͋�o�W[Z��mj�Vx��9�n�[t�5))�5�--'?���H��w�Afo �U�����t4�l�G?f)�2��_o	&�rUn��=�M��W�/K͏���7�G%�;��n5 �q���b�2\�����`�uj�Fw����X��3�v�,�Luf�#i)�߅��MXC��*�6
e��}��5�)���$��~��V��uu��_&�Tp��BX���Z��X$���c�,�
{D�v�/���x�Q7�������i5�5�Qk��s�1�|�R�}�(��'��{L�>��&R�?��t�59!nS�PA�2hH.y�G����~��Ȼ�=�x��,��n�\���S�����͋�2�`��W�2��n�b�g�)�T;9M�*��8��>|�mȶ`Ǳ+�	�V /�峅�M������;�ݗ�)"m�@�A�t����9��,{^�k'�C�L��R����2��p��G�h
���p�O�B�1��3A�t�yc����K�4�w�K�]�ߺ	c##qU�A���6��{CW�]"L���?N����+�z�(�K��XƩ���*Ԩ�L�A�EΤ0�a��涽S�cF�����|T���L��"��[�'F�~�8�ͣ��  Q���U�+?�"��+��<��q~�zvO�w�Ļ1D�j3�u�*mۦ��  hj�U8q�
�OE=X���Y��:���U���uK��_���)��ʷ��QL�P�&�g��24y���5^y�1�4�FHb΅�9t��)��PE)gt���>����e������*�g����Q�ya�=������JBU[B���h�"\ot� ������}�A�Z�U��5>?�=���z�)e�S�5�Y#��}������9ʑ��є-[�8��@U[�u$7��] �f3�HmA���X �=�(w�����:�f�"���@�a���M���N���G)���j2�<
�Du7:#t f��-�e�*9v�Ժ���M��\Gj�I.�:a}��o�9��J�#C
T��zF�e_<3�ԃ���MۻG�9��]MuXJ�p{\6��&g(u'�^��5�h�2[��X[M4+Z=�ߘ@������?ţxJ�Y�9���3?��X�w�i��3Ȭ��G�Bd$�F�<9�
d��Ӆ3 ��r}|:+Ii|�y��z�M�H;��5�̮�����{��R�6��7�n�>*/�i�s]S�����P�9�N���YY��w}~�2�r��:�
疮}B�tDPo�j�7<[���i�Lv�~_Њ��y'8W��tCGB����:w���o�����g,7�g���^@�~��I����V#�
� �_!�͟,�ta"]�,�g��f��wg��Z��]E~����-��L�_��K��]q���!>4����̣�,�2���Eۅ&�l���QLb�N�X���������$.~o����$�sWsl�ʾ�^�-��e����w�A�eR���Ⱦ��BFɕ)!��wf}�00��?7t��\���@���;�O'��K/m��	��b����~��ַ��3�����	�:�D"�y�Z��=�P7D�F�֮����W�R���f M$Kl�B�4˧�ٺ�Uzg|�1�u c�Z���=��6��E^��t0fέL�Mk�/�d��%Ր��,��Kh7��^"��\��c-��[��9��_��=Տ��˥�e>6}��$���ޟ:��B$5�Z��Lf��&g��!Oc�P�2�R��;?q)+&�u������z������j���� ��*�۝~�YH"�H��1}� <N�XA��B����*�T��36�#95��J���a��i��c���,W��D��sv�8�X4u��]��Z�pN�q.V㹕���B��3�z�GJ�@�N��l�P�_�1_iƺ l����
xT��$�ݢ����c��"��ܟ�\��Q*<�f�힯rO'�_)�MdCv'4׷��E2���]�ǷB]��CJ�5����"����ܘM=	5��\Y;���u�E	�/ĩ�@��$���| ��OLe��P�Dغ�v*k�߃��~�8������C�j���C��/Z�Hs�L����u6�r^���;W�1�]��
w�ޙ�4|�X�(3ذ!�7x�K����L�i�����w`�2)V��d���'*�]�`SOw16���w��w�[\H��n򼿏ي	ok/�zǃ b��'���G�iЋ���Rl�9�:�ܼ�F-�eqO���cD�����4/�������K�N�G���=�[�,��V������_j^�Crx�R��{�r�FY̥J,���H
�LOO�촬��!��V�m��=Ĥ��e����B� _�Wh0�G�S���]X���I2�;0�<��,Z&�ڏXߘ�<���1��yጊ�O�q�g%'!��R��Hp�H����1t���í�T�G���)�s1�ɔ�D��:*�^�H������І�5�Q&����=0Eہ�*�Ɣê�-4�ۧ���D(�����>�����JB�#͇4,��t+�A�o����ިw[T��&��y��18�V��g���t`�[]�
z7|~�"?X�m �����\���cp�Zڥ�;�7j�L��eu+4�"@FCOX�@�<ASj���p�~��OQ�D��tbw����<n���X*�~vV֡�8���U,Q������9���c��j����OS�.�oRU��M ,��U'��7�i�������^i�l��:y'�RH���M^� ��pţ�ፑt5LNZ9�S��5`j�k`�_x?���/�72ܱ�h���źTL�C/�T9����5G���lq3�ik�����{U�U'��Q���HGg�'7��X� y�R�.iޞ�$��|N�����C����ı1"���J=Zs��T�~.~|�fٽ��n�͗\p���R&U{��%"�w��wΞA67_�k�5��*v��g�dl�ح���tAH�L���r�+���������%�!7Y�1p��e�{2����6���9���_�ր�@�X���\��_w�9��oh��x񤒀@�)���p�m��,�#z+��5�ʷM9*35ۓ �C;T(���"K�S�gl�
�m9G��E`��	ە�����NK���(%<q���}��:�i�p=�a^�G�A;������$��R�FAC|�ƈ^
a2�\�	��<B�s�%_i���Ma�&��jW�Ԝ��Lh
8^��HϮǢ$�{�.�/�\#$��rF��
�;��s-t{6^�'�����Hi��E�P�}ņ�B�#� �C�Հk�.
��V�]�ILq�.�#"o��$e�_�����i��O{a#�0Kw����;�(v��b�%�f�܋l�Z���&,�Ͳ#*�%����V�]˳����mN��x�������0����<����3d�@����
�����Â��($�rGW�jyhf@m����X��@4�
��c�wӃ�os��/����@c�F7^�}w�ܜ������e<�:0)�W�@ڻ0L�G�� -�DzH�3���v��mo ���A丯8h�n)�`y�2���<`M{�v����%T8`�Ȩ˄&�.Px�*��mȃ0���a�S�����G�F�=��r;�|�9?�2�Cw�Cy�-5��rӌ�2DW�ڣ�ak��[)�G��� &*NHp��XqE��`WZߋR��a�) u<�3GQ+gͳ���e�脷�>������c�3;b��"�%B��LBUy��2�/�n;Ź�^V���ӑ��++	w�>�����SK�ƹ�~�R*��EOW�k�%;H���`ۆkT��&�(ʑ�l��80��T�XG�KY��4� ��m2u��j�y��T��E�	F����8+\���HsCk���Y�1���)��xz&0�d)E#|5X�z��F>+eP��5�7hQBVAœ��Ppbkf��&���C��r�S����*��4��4�|�R:IOp������UXQvپpl���p	N��i�Vk�t0���n�{���l�R�\�qh�m����<�1�לM"�d-�τ�^Wh;�����0�2Gű���yD'���R��?��čl��e�+�|�?�����bgo>J�'P��4D���2_���W�v+�h~��쩝���>�44TH_�B��R�k	���=c?��P�E(������h�@}�{��ձ94ҁ�hg���@(�=K�r��ԦW.��%*���PWCf��$�:�r�ɪ��t�	�U�8�q���V<������^u`n�H��CTb,�;���I�_��v�τ����C-`k���#4D4?��:̞n�+�k-��)1]�}�Ą��G��e��H��6�XDT 3�� 1-���+���3rV�VirG�ZO�H슫j���K�^}������#ҧ ���˿�g�h��/��A�'G_L{�5��
T�K	a�M�_��՜I������"M��_hL�q�50�^ 	x���<�aH�S�H�a/L��t��v*;��EdF͟�ɕ��m�b�A���]�3�Qy.�5��)[��#��48�$,d�L�<�B�\u�ƏnjW�Ṃȴ�jv�7Ȉ}%9���mc�5g�(L��<��&�N�Ѯ7�e��E��P�K�6��%����y�y1����n��F���,����QX�ͧ����9������f���VKӽzU��K|B�?g���KA�tr·$ B}���$�n����.r|5�n?DSg=>˯��p��L����$�p|3�B׏b�~�k�Ǥ�0��k�Kٰ��b�!Ɔc��.��-��T��(�vS*_ԯ�7��r�G�O�0�x�A��+s	�@�P7�0�m����.:U	6[
�(T�{O�M�������EZ�}Yu��T�o����WJ� m-���r�U�ɱ�IL�tվ�V���U��7Ͽ�3���I?	d]pu����,s= X檖�����d
��6R��ge�Gн��n�y2���)��A�l�LuITʃb��wX����ȄfQ�WZ��!��柚��O#ͯ��3��O���qg�~��n�m�G=7�U�<�rt�Խ|r��P�z�1�,����l��"ԸB8��A=�p˕1��O�qq��� ���4h�8l�uK�?6�^�'t|��+&�*I��Z�z�VYi1���"��z�R�C���<��]�y�-[�-i�L�Z�@���y�Z��=4��+�yazu����R�DV���f�q�b�ҟ��A����t�r����o��/]����-pb����ѭ��]n�=���ll��G��׳���A�j�R�fwX]SLO˞=�.I�M�V�+ �A���NH�]����=�����kV�;���C}����ilwj������������^��ǔz	]�������D����@��R��P���u ��T@8��o�0��Y�lժ �̉ya�-_�G�q�W�܃�w��P�3�p�v�0]V�J���T��K��N8�1���P��E���T�ktQ�X@"����s���������PQTlM;ˀ��B@��3VQ�凾pt[\%�>M��}3����Y�}�b0�/�z�Yy��&��b�zDZ���F*Ѵn�f=��ښZ�6K ����ա�0�Tt�8N)Oƛ�a㭥-��P�ܥ���;����!��k����*J��v-�\���K6��b�@+a#[�����eV�1&�����Mz̦������C���hX��G3@��Or��2��Z~u����2b����n� �һo��|*���?��#��������e���,�zg�S�=�C��9�����4D���o��$�GC�w�L�I���� 0$�$���� ֱ��䃚D�u�^�����Fs���7?&�����,瓐#��Ii'��ۊa�5���E����L/���Ϭ���S:xm<�Ծ�e�w�n�I���=�����.^��&��G-Y��pS�`
fb�H�N�fm��$�m����xY�F!�����쌿܏�F�M���Ȃ�)��[\��ר`��u��;�+AUe�]�3�s�2�W�|�ΎΛ
Ⱥo�Q	~d�ؒ������'��v�U`x��0�Y�xȄ��g�����+�P�_��"�Z�c��}��@y,@���+��-J��1"���^�������+J�v�wȆ��џ�c���k^����K.��> �hh�gS"��F��U�S�*3�M����/������b�;&�H�]%�*@i�!&��LJR�C�� =Ӻ�b�6:g�c��1{q)�t�f� ���+�u�OAn�G��~_,�lA��r���R���k�F�)aa����3pp0FsvX��T�5���������5h�O������V�³��*�8T�����g�6��Xཀྵ�IP ���_�1��jU���K��v��l#I��0=~��Xxk�P=��+�/GUM��!�5��6��(�ج.w����Йt��1�H�=�+	���G��R�r��R�Ysj�j�~��d�V�GM��*��LD��v�7��-¸h5
�pE�Y���$Ѹ��t��k�R�9�Zu�3$�s�q�����IgQe��*r����@�����P�v�J� ���5���D�s���0WG�:ڒ��+�5N�cX?��U��vg���mxq?\c~u�"�e�PeZ���!��j ���)��Ù�ke�U��͠X*�]�N}�:l߆�d�%��P���1����
R���#/*P���%�?v{��;+���z�78:�!8�����n@�y�a��D���V6;��F�@O���(�l4/d�;���U��Qou*��|��i]����q�?)t�+��������~0]���Aփ��N[��=q�[Q����9u�e�C�`)D^���-�Vk��8p�>/���e���u��}�߳�O��#'x��M�]�X*"?�X��#9_x��F��?�Q�!(Z�[��7c�B���]g�̨�1�ٟs�*K/:�"i�7<7<�@�>��=ar�>��/�cٓ6�+�7¯����yw��c��^�s�쇬�|�N�N� \'�0^6�F�j�\�g;&PDr�`�v�r��9��i��ᒨ��s�����N�MΟ�O���7)+j���>70��^ZNf����3k�~ʧ<� on�(�6�X������ A�:�l7�A/��g�2sQ}Y�U�с2�����9R`F�ú�-�(�3!��LJ�i�v���U*皡�њ����/�?�88V]��ʍh�QԦ8bi�)�lx7�뙯�e�:���,��CJ�Q6�vw��G-��j@{?*y�܂*�ơ�4�t@��ϴp=_Ds�㨪'����	.��,���$'b������KFИq�/����a#ջ�jnuw##���խ��3BR\ D�+,�&՘�!C���kf��Av���Z����O�k`�`�x�+�6���B#���6��;B;[h^�����ݢ��M��kA��]��)�!�+��m�n����{���PT��d� �z=��k?��/��s����W��b^��X��9�κ�:ݏ�(�3� ��XJƌ8�K�U�hn/)?�22	��?���A?��L�i�y��C��()����s ���t}X��)G�v��{��~�@ŧ���.�z�������IGW�䒮�!�d���1S�tF����{�<2$��������`�k���cE��p�(��=�_�"9���e��m��.�N�U9yƌT43�=r�~�aG_\c �}��.9�����cC�$M��VQ_i�%�+�u��ʠˣ)N^ߩ����Zn�U��[fE���d�r�����B��Z��PD�A`�R�D�O1��y���}����~�Ψ!�I�^���fLE5�M�@���8M��ڑ�vT���8�?��ƭ�pN��~�a�wIn���,N��P�Εs���N�,��7�֑��z.�p"=���r���r�q%�u�짰N�l���2ֵ蚻,��zu�f4�����eFX����I ��.s^N,@��}��`��˸[��k�>0�y|4��ZZ?�j�r�v����!���3�6��\�����7Z�������Ne�/�z��;�RT�R��Ҕj�7����븮}%;��x��?�z1�\�?)� {�-���>�ӓEX�?B�'2�<���﯇�l�f��,dy�x�q�[c,FWB�6*�$��X5�Lv�l���� V_ڗ���曶&��Ht���G���a���bNf`<˅�U����*c���<2-7�P�ҫ��� �'5"�CJ��+aPfҔ���F�̺���,=�c'�T{�"9s�^5(O��v�����E�:5g��۬2:ۿ�W���Ʀ�%'�;����8�T�;�I�f����wF�Թ����ݾ�^Omn�g}�L�L��ވ�k�ٓr�1��z�0��܁��H\�0~�h�{��c~�j�#����4(���bƕ���N�O6Ξcc�W�@�fR>R7��E��с���r�؎^^�@����Q��a���AN��=6�x n.��sLM�5NVH�G?�����L��.~̌#��d���AGٴФ�!f�7���>B��^����oya6�6(f�p���!���Y)������]PM;t�(�4�!^
�b���$��ԗ��O��ۈ8,�)$?�M仺�?�w<��++������P_���Էգ*����is���n���r[qy�Y���˫��:B��
R��z��2�&m�oES�V�"�J����켎�����=Z�Aj�b�:�ޢj��5�C�
t�d:^z7�L�r��?z!�
�M�ē�H����`�Q��t���H��^~P����$H"ˣ�e����E�PU��sәROJP�ㄻ}@1�+9&��3(*�؅�U7���-[�nj����x�ho�������>�|z����ɒ��e��R,
��3���'q�~H����{��(( N��]�	�^��R�
�%���"�R��"B��C��n�D챭O�:T�D^̖�|�I1U5��\�H-��7�|�k�"���|������.��8��-�6��J��D��k��?��	��]#;u�iD&�Z�u�v���d"�i�>,��}���pw-�3���M5���Ar�"ӑ��J}��`�l8��R��PF�#j�w���1�	��ً=��	�6Af����=��ǃ���E�݊H59X��Z}@,л�Rx$��3�7�c�'̼�g�}��Q����Go1 ���G��^��HmC}�Z	����鞿$��#�0~��Y\�,�_M��b�p�&�F9��"���6̓\��m�����tCF��).f�����P(��^���<�u萦x�m�ٺLNMg䋍��j7�l� [�4��(EQp*�v��Pd�������8�0ɉ^vxbf�F|�<���h9KGV"$	y�� ��4W0��s6���k)/�y@�\`J�IY��e�/!��� 8Z`)PEA�q�����?�v=�)���������2;��G�T޻�.��C�ܹ:�#�jG�1����c�dz��	Mx�&�M5A"lg��/V��>�����M��PT��V'��I�r���J|��E��@��a������o�G�j�_��aYУ)9l_W�T0��{I.v5��D���(�Y���TП:m�9x�D�C�õe��ws������ �;_�׿�����z�% `����2���۵bf3�1�򁽳5cR����oBv(�&߿���-�ϻ0=�ݹ���	%Bx�sY>>W4�l��\�gM������d8�ˠ�b!��m��h�@�i�����e��p����rb@�r��GX�D �Q��Q����d%o4k�U��~�./�*C��5ai�� H��s$�Sr��5�_g`q�����XJ3u�}cd�lt�0{�����T�R[GW����������l���(l�u���w���Yn�6�ĩ�F(g:�Q2��)$9�� E���ˋ�;�r��f�ؤ;��U��˻�tj��*������5�Z�d���R!��?w�=k�V��
��;aiH<�`� �#��@H������I�F
�)E!�#��x�a|�t���L� kk����~���j�<n�n�����(}o-g R>��})�L�D�I~������U�K����U���W�';���ݼQV�:D�H����<wQ��,JnPB�s���YV�ı-ne�C��vg�X�7�9l���2K0aL��
�H�Z"_3��[U]B(�N>zW�_��Z��h��Ak�0r�?���ۉ��c����l|hi$>P^��j�����+�#1�c1�\�6�h�TlB���ԙ��E���. |􈜼�M�k����+�.�_�b���˝�#<����U,l^LEB[s�>�����'�Z�ϛ[���R���2W���R�Zl��%����G������)�<^[.���kQ7#�7����sO��0��J���b�?���er����D0�2���K��%ֹ8X�2�Q��[�>8�i�!#<������-��]��92��9��Ī�0�͗���8�N����:q���Rr{��w�	\�䋟;�Γ �Tl���4_�[��]����WM�]6��s*��-+�^P ja�=*�ݍ�R)�Mh��G{Y�%�e�.;Մ!�,��j��E�L���Ϡ
x�4~�ņ���UN��׋������H)��l������SN3'l��T�D�;�Cz�9�( ��hZ�
���<���"]`h��:�ӧl9א{�)?f��L�R_�"M�I/{_����`L0�Y�q�QiN5�����<TM�s�V#_�R�o����[���)Y��ą��ܡ�;%�i&�6��3R�t�E1�n�I�g���^�G˿�wޗ����p�ð���-|�ǀȓ����E��[�i�UH���,�h?3�z��udJ��Su��F=�cp"r�4�u��mF[mڊ,?�����x����?"��n�Z�s�s���!��/��R�08݀2UC��]'����F~h�B�<j�y�BE�'��(9�g	���j��yX~Ka�p�H��T_���-���]��§��R/Q̂q�PZ�v�q��x?H�v��ϥ>5��g����������iw%r5T����?\8Gz�Z"i���v������#`b�6���������G�o�l�Ȏs[M1���Ѥ:�E�`p�M����W;{!8��d�A#Щ�`D���UP4"���W����|6巙���#n�)ά��f��l���0`Y����Ϗ��{VD;7rr��r=O~�0X�Y�B��&"��0�[-V�i�`�m�c�Y:���%����� ��`�����Z�Z�Y��濶�}5{�r�{1�ų�%SB��j>�R���&�VӜ��0��]Cn� |�R?k�^����6 劀�]1/䭎�vl�0��73�a'G�:�.2�Ui��:fвW�X��hC�΀N��]WO����}xi�h���S�F�"得�\6M�y��~0������Nz�ļ�����Ǯ���R�6PZ�:�},��}UY/�dV xͣ~ѓP�TGO���<Ǡ;a����"�i�k���z�W`�b=:����3BP�~j$���c���x�B�z����dW��#�'Gc�������}��)Bo������D��CN���>�5���q4�����[�	��e�9�#�|.���W�6�֕��,���{abi/6o��\�{h�$�ħF!߳�<����v����y���5pP��~���rQϜ���1)��C��g����w�>��1Nn\��σ��Uw�l�J�RU�D�ݼg�2a�2kh3S��a��='���&���³�>�(�+�qF
���VY�u�]�/<"���M�χ��Q3�[��\�<�*��.�Bx�a=7�Pǣ{8k�����]��&5��b8��G���:@�@ �'3}H1�_Ps��PX�=[)�ŷt?�#�.}�::��J2�r�/����#m�9�$�����m��)����*[��b�;eS�j㴝�0\x8p<%��rPN���4�ԛ�ӭ/
n>�1��[}�\�Ï�jf�2�������U��͛��zi���^g�+�Kt�t�F�xq�����n�ˌ��VY�V����ZӁ��	�.T�Z6&d~$��1X�A­̱'GWLT�P��8Y��*l��7_4}�4��������1�Q���LyEob�CC���������y6�kP��=׽��9lh�߆x>Zv 7�"�%�B���C���5sQl�Ұ�h�O�"����ƭ�h
�,G���e)�i�kYϛ�s�&?���t�Z�ǫ7��+�!�*�݀����m�Vp?4Ą�(!��7���T������U쥙���eլ�c�T���Ub*(���.�t9��8^��1h�'P�Ge��������Hy}O�h3B�'Ыyzq��(t�(���!U��k�u��An��/L1�Cچ]	�N\-���ʐ�(�g��:�/��ΑN���&SK���g�K�ڌ��r�����Iu���g��%���w�?$�_�ԉ�#��As�ܣp[5&�Ko��`�ϜHJ~����L���o��$n`��M5ӺTW�kƑT1w;��U��Z��$�Eل�Ի��3���\D�=�^�I0���ķEaV�VFy��������bA8��p,���� q����B_O����<6��Fx���<���P�Qު7� ����l�I�s}��^p!_I���	4��S��Δ��*'�:�wة�xz�a��I=�P@bݘWyW�ƒ"9
hة
i]�pܤ#��� ��x)�M��Ô̉��|+mw�����uN)���(L  ��Iqٯ�^�? ��mW2]!�"���2*� I��!�)�y�=�-�̌�Nt��YN�����nb�D԰ⷁ��Ц��4�2D��E�aA�����ȭ���p��#�\?QD+��װ+Ō��ɚW�%�{@a%�,�*���B��o�Z�t�5;�ӡ�h���XE�S:US��E՗�(N;���\�q���� (�0\������S�u"���|~�-Z�NS}�T#H{ 7{-.��|Ck��)�R+�M�0S27EO_}jb}��=�C��l��)��8 ��N���iajțu�<� ������, m�%�I$���teƁj��㡵}7uz����{��k	%�H֛�Ʊ���8ua�=��n��
�AU~�`(�U{��9z�m��?�$-6�<�E�o���dg9N$<�F�;�K��2aw����ƨ�z�A��Jw<YżNt��vB�������D"u�J`����n��"�ەs0a�S��wS�9�yi�)�7�a��h���f&��	6{�ɽ��T���!:��A�V�iA	GMJ� g�{ss�m�,K�
�槷t".W���e��BE�q8����@p<���8s���ۻrR	yx�����W�'S�!	��$I�u�5�!��3�o���7 ��������D��bߵ$?{�"N�V��7~�YB2nv�+�Riɯ8��չ�ud�
����̻���I�y��CDQi6���c��_}� RO��4�FliѤ�ꎵ�J�v��-V�w
zCׅè�֊���өy������Ё4
���Db{�R&�ș�]�~�t��u���5������05Ѧgd߃�C8�\g#���M,_'3yY��
�"Y4$�O��3���m룲�!j{��;w>0?�����7�&�SC7�^���ͣ~^i���Z9v������0oo�,��n*�7I$��z!���t�ec[�(1�Ih��BSV�zr�s��E�:�X��ND��q��S*E4�Ǆ�3$GMA5&��&�M����t�l�gE����à�X�)��,�뻿�]����S<�Iܕ��p|%R����Hh�6c��0q�Da���K�J>�Ս����X�i����%3���Av�2C��z��ә�~T������T�Md3���&qU%1YUS4޵KZ7���%s�ThK#Z�[�DR:��N�j�Z�;~�Ⱥ���S�DE&�����*�3=�0$}�F3����n�ּ�w2=4�h�=�PŜK��u�J�ݧ��[��@V�U��N-,��j)I�F7�BE�_��ӚU��X�DP�>��ay�o��Gl�GU�1�퐾u�Ҿ׌��5�������Bw��8����3���������Ԥ�I�#�:���F�%D�}M���ӻQ^�h�W`K�=��1	��Sz集؍�� ���E���A�N��*��(�eR{Tw��7w5D\�͹N [�������+�t���~x�OOC��o�%z҅η�d�V��*=�K���t!������A	x��8r�T��:9�)�+@���"���k��"�eC��VT��7u��q�׺3���6(C�����z����7�h��u�&w���T�J�g�w�y�m�mt� yQŠB#�9¾[�oa�r�.DR�?���}KXXvě��.ʹLr�D8�,i>Ue ѡ���ʪ�V{�Ùr+�����H�R�ɻ���SF# J-�(���=�����jA ���&k��BK'��.9���6L�8�Z+��'yz�y$�H��l��g%e�DĠ���e�S��ˊ{���;e����6��ZU�����b,�������J>����C�,5tH$�詳ɕǗ��~�Z�S�����$-�1�H?�a#c��H��z���J�+�K�����B܍���4)1�H}���U�]�P��{B�����q�����ʛMa�6;%���":��E4B�fqs!9@��3���JK����@�ds�M��"<���'�Aݮ��N�25j��\8��&�C1	��0KZo��Y�d�b3р[����2�1�D'Wi�r�w�ƌ|t�ǯҦQa����bb�Y�/j,2P%=��9~� u;�Y9]~��V�}I8b��k����P�V���t�,�c�S�|������Xr�g0�����7���s�H,㖇@�bUF�phC�:_�
[!�fT�1��=�Ʒ��6�[��g�3O)��]��yֳ��&�'r	��9�dZr\K?����U��K�w!�eƳ��@�����}Ƿװ�Q��IA+�������T�;��� �@@�3c����ݩ��5�cu(_גH*��z;�LI
[�V&�4,F���O�>aN$d�c�i�LY=־1�;^/����&GĞ��fh��KQ���ͱ���`E{Dږ_��?�׺�.�|b�p�w�[��̂��2w#�ʞ4�BIS�ZA &	�ұa�KkBS�Tm2���}C��f{qOo�j1��j�y�[p�����&ʕ�)�
��ebfӻzq���ޑw��^�[�)F��� ~�(�/���9�)��\u*���ԍ���-�	�A��8�/� 
�ڣ�Bf�`���ׁ��P6�$��
�G�p�@��v�\BEɣ���!X"p�Inb:�=�B�����@ѴR��Iiu gmW�$��R��Ź��/n��I��r��Gϐ��[�Ъ d�E�FԞ�.!��3�r5��eF�g�:l �LA��LVZ;
��`��jJ��O�ZF��B >��s1txL��{~�����l�%��w���!o�) /�צP�Nu�S��T�1�t� 0c�J:xR)#U�A9�fB�S��JMG������/fO}@�/���Z%��c�� ��W#f�~-��o���I���i�]Tdn+u�Ke�,��]䨮�N|$���Í�߹�R��)�Z�d��H�U	҅==�'�u�,�b�����N�,ˈ�;e��
ca7ͪs���!e9��j�å�fs��)�}���/��6$�S����I2�B�g��F�wz��=���,�s����u�w�(�]=��6���@}hŢz:�a.H�C��,"�
��������믾<�3�Al��uu8ǡ�F�c��%:A�u���C�x�K�nT7}�����'�e��W��j���uH������/U�d� 6U��OAj�1ܭSOs���[�ob��
�PlDJ���)k�^C�lD�S�}�NJ;�c�;8��Ĺh���#��!���	�ivBߵ�ޑf�![�FMU�U0�(w�u�}ʦ Y��^p���MN�K��%'����P{iF��w����r��j���j�[(>˂�v��!���́�4nk����Y�$;Hs�����f�LA�H��(7��3����D*��/2��3�j�W�|"�`��a�[J��2e��ZL�]�SS�?�02�,HE����=��q$:���G��"���005r�X�`�1�V$�{Hz�Rـ��0�۷�=J�{˩��~���d�x�'-V�lA9%iH\++��x�G3l���)�ďT���l�YiIE��9�z�|�K���I�v�s���6����\z���%r\Sa�gE�l�v����O5��"�\@@�{�Ss���#��}��QR�!M�I�r�k���Q�,؉ x���jvs\�TD�C�2עϝ�tZ\8C�y������[a�B:��b��a�ì���iyy$D�O�ݲ���[���
V�Ђ���b�5�3�dAa��hrY]�:��yH9K�k�ڵ'w��P(̩-w�Z�)jx��ﻨ<M����~�u��!|}DRV ����I��RX|�އJ|��bĀY� ƌ-�1�J��_U���Ys��bz|��)�T���e��kv��hD7�i�ۉ�Q�Xh" vKT��1[.�x��+�U�¹z�!���T���XM��aq`ыw���UZRrNaLv�5Ӽ:�2�.ՠ;l^v�V��7Ơ���si�27S2�����#M�t�f��D��d��İ06%�͂)К���4=c�4�,OȠ���,�ZX�X��
=n��Y1��9�$vK b�[�u^��-;��>ý�ݍ����w2�1���"Z�#"��FzS��\	��'G�lH���rY^��{�l4*������k>{:�ם=����10xJ{c�M��h�	��m�2h�xF�)�E��9�;�[����:�4��7f�تd�>�M*����ԙ�vd۶K����W�^˟�7��k��cRp�vV55���o���{O�w.���u;�߆	.'�%s?��n�lY��<�e�s��Ȗ�c�cVz���ay���¦ƞ	�fN��M}�ak!��&
X�h�J���N����~%�Z)����!-\��qd͜H<�n�-�]1��\�b�T�/�F.�K.���?_�gG`Ry~_%���K���{QX7+	w��:��\���7w�Q��i�����dU�빾sD�"�y���N�w��fϚ-P���A\�5L�Q~�ga���fg��..vbV�̑��ؔ�[[�G��y68�{<I92�!(��ؾ�zC�]��d������d���M��㹱�B��n��5>Gov��l�����-akN���o��zƗ�)�s�3�0��v����(V���a�V��F� g7�7���Y2ړ�@E�r�����[��8��฽u�J89�d�ix� M�sU)��N�e�4�FrAb�+F���q����٬��l}D������9�[a9bB]9/�\R4^^��1Y@3��+�4�\�{J->����#^x���-�c1��~��t-�K��%����c�M��G�2r�_M#���kQ��դ���C�%�b��;��%�:?7���&���߬rO�X�S��5�V �CR몺a^,�������X}��ʖ�(�.XA���|�>��@�!俙4��d�PzH���PL���{uz�A�����o�`�u}�
u��EHH�?�Pl��Ӟ�`���ʧuP����XL��P��|;C���T�q�+�X��e������`�lˮ��;������y�.�󴼣%������C���y���E��2���hq�6�L���������6�-n�;�k�X���Y���
%���
4;I\��٠w��J�KT����w�31Ig�3 �<��dV���=��Տ
��Ԣ�!sϊ��(|�.��Ø~k[A�	p�z8Z���Y�E���s���qrݑ���c�p���X��#�^x�|��n��=2�l?hR���k�$�dy7�>H/�, �ly���}"�0�^�����k
�$tWƚ��O��^:s�}I���CE`�{]�uo GD�]WF7t
w�M�@�R�)n��5��湾ב"*��gX��Q�����<��,���x��;b����_���Ļw���O�;���3��F��`uH��YZ;�0����vK�C������_Y���ڥ]��� �P8I"[9����'#hH�OG��p���ťĖ�=���
��F������[h����c���܃L�T�ԍ( �c�L?5DY5�>��k��:���:�ψ'9Ƹ(G8�5Θ�U��٠�#�B�-��kT�)���V��?�+ِ��H��<4��6��&�ލ6$;h	`��QҦ,�2�`Ԋ7�
��X������4\oK��)��8��M+���Q8N��=�ڏ�d�.��bU�t�Z`S���ARec.z�@+�Z	Ro��˄�;o= ��ͯ���q���h�_�$T|���l��$"�J�8�2�����)��Lg�DㇰxtQv+��C����B$c�іQ%�E��l���d�X�wx|S��|5���V��^��.y�4���?FK%է�jq�"���uB_�A@�{{q�� _@a�+�	��JeGUT6O���������I`�a�\2�h����FAa��;_��Lx�'H����.x�1I�������ݠ*f�-S4fҀ�I!23���� �=��kK��D�)K��*EzBR��F�Ҵ-k�Æ�q�F�:�^3�]�:*�^ɽ�T�.j:���W/����F{�:�e&��)�rQ��/��|a�TW�_p���3����p����@������Б=�KOF�=E� "v��v9�閭�ܹ�nJ�����c��|7L��^��鶏�o��H�	|��V��!�\�^��Fg|�i�� ���W����,7�˓+�d'�5}k�SRn�s�L���	0r���[�����'E�h���?�_�7#bvb�r��v�(�|�%@���C�����d� ��.N�f�jHi#d#ό���ۓ@ �:q
fX�ͱ��ŕpiB��%����w��%�IL�K#,��=��0�[7�]����d�Vt7�y��j��~������Gqd��q7�!d�j�f�@���B��I��"a�9��:�Y.tH?�M"�&�~�C_i˹۩�cG��R�E�+�Ί3h�Y}k���PLkVohzU�C�d��R�>��0�'���l7Lr���Ab[��=tϥm�^���0���qz�a�mk�'�T�63�	gcC���v
t�:G0K5]��D,L�����m�+I���sY�㍂�/��c��B!��"zp����j����]���¯��/!ɷ�S@��{������\��k�G4Ԟ�M�\\�2���25��|<Q,P�T�(�$��t����')@�@�zc������V�'�rtv%���� 'Fi��u�����̩�Q5�OXE��}/*�u�;�`�O_}�O����Q�cG���>)�J��\H*y�l�ᔷ�U΂D�=�#+;[�,پ�(��N��q=)�&g�~/#f��-uOBZN�yiK^C�xh�7��Kg��xl�⣱
�7�fs8�Y���5�[��LZ2
*󌪡���fȎ^^R
�6e ,��t�@(;��KP����q���� oʯ�UD�
G`) ����1�Jq�v�)Bq��b��8Tp!�DH�����q�ڴ�TT���W��X��G��v��I
��[Pf_�y�X�l�ډgAM�h�ǀ��*���<R���x�g��Ց��"� ��ܐ�"ˆ�h�XJ���,�guJHdy���Z��'y��w�rԉ�(ڿ�9�W)���̱�0/�U����Zd$���$�ʶ�
D�x�!����j��N �]}5�	�Q)�S���8zd9�x D��ѯ&&ߺ}��M��u��R��%M���4��ց�lM��r�s�B�iՊM*����.Va��=��F����?�9n�����#%Z��1��I���Y��T��DcP7*�brp��%w����*�Z����j�ϯ�f�΃L��Kj��8^�P+&��@����[ba[��d�h֕����4��1����4�FS��W���[����ng��Bۃ.�-��d}��δ�>�{x#��S2�����b����h{ƫږ�L�o�-#ur��}��\��h"���2M����*�u�t)�(nA�_Z+C��e��^�l����̹Qch����d�j�C�01xԿ���N�J��|%��|�Ө҇��#����x�1t`���a�ג\�q�CH1�[K�J �����:��(�({��� {���ܪ���2%����%�L�=! �@������ �Ξ�KJ�9��cnP������GH���mZ^٣�&��'=�Cd˳�#�p���o�ʽ��4� ]/����#�u�zݛ��s+�x�ʊ�s���_S̩w�t`6T�ɂ����C�F�
�[C�I��O�С�B������
���&+9����ot�X#�4tpVh�W���w��&���%�^~C/q�y͗(��!fO�|��8��&$�x�}4L"���lJo��$[�k���X���oH4���",��I�Qm{�1��?rXM^3 �0�d�4~���Z��pF��_g��s�[dǼ;h�9�6\?0;���i��>'&�ð������+NPί=��F
�^�7=���\��1�j���q�世�,���x�K&����_F�J%�1%�~Y�'_����-�n�
�|���e�����]��ݱ�^�k;�#�pAA�B�M�����
EŢ���������|�@|?��)�	j�!`���ð}+�m��A'��#v]Id�Z���}�/Z]�Sn�_�������i��m6{;�i���������W��w�0ԥK��!�Z��*z��