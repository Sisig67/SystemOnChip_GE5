��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%����:P�f%��mnn��Dm�n%N�w
�cM����_�WJ������Y�G%Ih��|�N�^��dTCȮ�� ���e�<���&���^P����0ST\�zn�6C$yV�4�|��*��b/w^?�?a�f2> 8���X/��v�W��'��
�uB<h���_�̻rxi��+(2��٦�����}�xcm�F�H{�����V*N	�� X?;�.��n�iKܼDd`{F�����s�R|%?�d�ڒڕ�إkAc� y��ŰXY�{�ZdhL�+�wա[c'�b����h������4ű�����6���>0Q�/$��Rs�?,F�Q��g��p�$z6�/U�OÅ�9��L���r+v�#���j5K ޸��X�����`�3��ﭔ��qbR�H��/X�*���CZ�-��zr��jD�b��RZ�/��%+��'G�o֦�#�gG�8L0iy�c�>�A��'���(���wz~�sh
�i��4H9+̰��p�r���R�ysڛ�u�������bŧ��۹b���Zex��{�U}\e�v�~�I���ӝfd�bR�$,s9^�G�ĕh�����eo,!dLYn]#��+o��ې̗o��uW�A�M+�a�M�R~`���Ջ�
˓��C�r���h�IKD�^-�i��r�4�Q�uyH1\5�ӹ�l<�9�3V�3�`�4���:g�q���������`�r�l>����2Hh��xC�Ʌ�)~$:C��aA_UV0J��2c]NM�?]��y۪�q�B�U��i��'lq�I���y)T15 QjDF��6�'5���v�h��5��� ������Oq�柑��{oETxIֵn�r7��_W����8�j�=,Np����M�2v+�_�À��Jf't�{��W�@\8���`jqQ��~铒(_XEV{����H4��wm�!IZ���A@�����u.ebO��(+j^74ޠQu��2� jq]��SɫK9[,��<�4��<���3��8@���ީm���6���/�s@ռ�x�[a]	AD1�"����)����4�>=C��y�׫��3&tU���v���c
R��&bVh��h��`c0�<���Z��~�Z���}�b�pr4��'�i�k녛g[>_��P�ߥ��А2P�u��RV��ߍ��}��������۹lU�(���d���|&���aU�@땸�Z���~g�фa��G���}��&�m]ZW�{|O8y99�
��?����!�九�!Dt����xN�f� e�.P4f�D`������fGc�z��kXm<ߧS
ʵ��7�򭿜�I�x�";��M�N�uP䤛4I�؅�[�`5ã�ջw7/_B5�����%=��r���;��ǫzG�I>ś��Avx`�L��OEK�3K���T�ѱ'~APbEւ��Sq��A�����������@��=쨭���gg�c���0�����~u�J�A�aem�o��VTƗ�.HD�Y
"$`.f�H�I�̺`5c�$Yn���q[��]"�f|�kn��!%R8+�G�a�����W��v.�o;W����n�v��'u��y���E}ŏҹ�����ʭ�z�':ꢿ���$(�9�r}6z@Wȕ��|t�kF������Z��=q��q���V��JBo����ve}{��9�>����T�A��EJ�Y�9A`�睕5�)	��p��������4�J�O
Y�Ң���%����eR��[��ʜ��l��{n�<�l�6�i�z���%���1���+�#��5H$�0毠�t����/�� �ʅ��*m�Ph~_f��<:8%l?�[����mG죎�Q�o���Uכ��\=d����(࠽m9������b3�m���/;@���qt/1�K�y�����PJ��td�n<? @El�z]\�W�A?�͡r�?ϗȩmts�{E�)��B�h����a�����T)Y"ʬP�2��Ǻy��Zͧ8�j-PlDg4�[r��ge�`��� oC`���j��{�R渺%*s�k���Po��-�MhE��F����k��\���V��#���?]�$(k	�L�Ͻ����¬X�����̲LC�^sW������M'��q݀wIF9�1�[�,�Fb���ajw�
��s�y+� )"�����N����Fj��zG���y�!pl��x�Mzc��L��6��ԣ�6�)y�9�[��qGM�����`U\�c|S�H6���`d�{}w	z�Q'��J:�
>&2rR�)&�<�x�$G��ϩ��垏��j�`8�<��� ��{�(�ª
K='�=<���cw�`n��6R�G�]����s~�_��	���ERw�a�p���V���w��6;1�ц������7^�Y������'���?��FZ6��_�p�����a���E��3QJr�+�~)��];��2{�ᚙ*�c�Y�B�I矤��~�9�ӿ@s{�-I�"�ϴ�����MF4�/��xc�^hL��RB��:'�W&��X=�1-�\�3/G���qU�d#Ƽ��G��;-h~y�6O�Ǚ��7��K=ɕ7ؼRT�r�7"B�䈔7�8��R��]����{:���^�_U�w���"BK{h�i(�
r܂��Dw���\����3D
�%�w�ϥ=l�}��˚s��_�i{�Β�ikq�.-}ؗ�C�#�b�!%2����P�cQϼȚ��I��9Q}K���~�4�_��Z�]�W���`�7Gؔ��x�y���q�$9���8��4/��j�&!�p�-��:%}5�R�T��'����T���R�k�?����@�+�Ob�����Jx(:悌��.��̦�%�Mh�v���i�'s���{1y2�E6(˽�Z��WS ��	H*%u��O!N!�Z���1=��U/��Q���2���1v�S��S��=�n�������5<&ټ��\�S��#O�^�Q��/I"�r�G
�}:-y��L���(2��ʭ�K���'W�7��f����1�5R�e�Oj��ͷ�8w��࿰L�?>�t��L6�6񄰘��!V��br�|��}h粚�>��΃�Jg�=��P�T	����ȷȖ�>]L]�g5��iogr���L�3V.��=i'=k�����*��難#R�g�$����4)(8bJ���P4
	ݬ|qAL��?����Ɛ(����/�^�y���߳��>�ֳ�Vk��&ܰhW���"[<�P�#���>�=A��r�����JDMfs}l��M�"0�]���Zz�+7>��y^Z��D+��/m��Hc���4^�T:��8�a��j�'�9�l�7E��c��B��� ��Q�2�p�!��n��	4�_����'X����G�^`��s���C��	���h=��5W��5S#��_r:��- O�h�A��+�)�\��xm.<-�o�e�MWvy�1���Ña�JȲ*�������o�*5��Ǳ4�����>�k	iْ`g�(�qocr�"WO���+\}P���ňa��c5b�΁��ꪶ�������K??�L�H�K�ԩU{��zv��N����sP',���g7�LW.JE�x�O�1Lڑ��)��$A��%���-e��dt���P4(&��cGzHM�Q+x
/��o��oz��]�}/q"O�Ϭ-�[�y��*���{"{V�+3DU�@J`����c�t���H�W}�@��I�<��t{:�yޔO��Gy��;k���j�؁0��O�<���Z �r�@	6֪5��m�1��q{�>���x�E��"�`=��C&?�x�`H��;�'�Z����w��%��Y�~�vn�|Q�?�)qܳ]H6o~�v/�Nhu�16<��Y^뻡�?��iw>�!C>�hP�wU&^��p�:	"R�Q���B�;rcq?�1_���|)�IY��im�Y�㌱6�]//��]��i߅ۼ�:���c����:6��U"� .�e�ot���3,�v^�_G��^.�,�E/���"��e@�+G�}��׀^�����Q�4���<�z��d�|�J���W��J�)6,[���r�J0��$���c�Ȇ����ه5�T�ԣA���jj�!��k�;�bR3���d"0�F9v����M^�L�6�nn���ң�ǁ�7wC:��%l�����D�A�f��i[,�Ó�2����E������P���R}��8�.���<2�ΫP��
E��\�3R��oÍ���ސ�V���M�>�$������e48c��T�����0`j�j�gX�eG�����w4����:k~IB�I�����>ki��]O?d�72qg����Yq�Ea�㻐��0@<���Rr�ٵEJ2N[�!ۻ;��9�q�!�^�r1T�kv&��7��bO�:�O�=KQ�~����	�g]&B�����H�"P��k� �1?9�����ͮ �]�a湕����@��>.�m�J;�2R��į8��n�I�W���ݷ�*v��a���-oy�t�߫^'v*��:�z <��s�O(��7�%��Z%�`��8��@��JO���N�$\�h#������n��������P��k��"`�z���GoU�L̀�8v+�R)�c[��&�SvL�f�\,}��2K�Cd_R��h<CY��x;��c�����G=v�@�W
4u��a��'��qf�ý��=j�¼�}���az�B�E�Vq�����F+��;����Dن�K0�!�T��ı����V��ί��h40��+�[_&�C$�;�,6l;j��L�vi��nV�>��7Cj��] �GS��F��"иKQ��Q��8�PģzE&Mnfŵ4��e%А�$�MKCUá����#|��U^�;�'�&�Ĺ�����p��V~��٨X8`�W�7�iE��t����d��_�Ԁ�6�#�[����75�:B�kb���qB)^^��yR����q2����=�]�9q䦯SŶ���fARM��>'�`�;�̣�����1i�zG�m�͂��5�& a����t��W����Ŀ��zJ�������r�=�S�|��(�f�^�m%ê����@CA�Z��i熻���H-yNS�6 �ʲ}@�i��Kv�E=����a�K�u^((�!�L� o�^r�h!~���Ε��=iJ{��8V\�<)Ř���(t9%�q��lQ��0iP`��x�X����S�Ų�chL:D�{�K���Cm��Eed�����U���� @.j�u0�k�)�b�,VHT�݌��쑸��sI�`o�)�_���e���3�4���9j�+B�Ngݯ; I���Є%̶�0���������Kb���:��-x��,�>����������jI�SD�kJ[��5賞g���w��`�!�e��a`�\m|�����*S�G������ȴ�C��0;!\����I믂a�+os��T�o=s�,+�>zb�z���L��#�޾�y��A��Y^^s���;R�pϨX��I�6k�/�����g�d�<�����?AG�P��uvd�rVΐ�n8$��B�f>;v�V3H�  C��D��~��5 ,d)�G�,C�~���{'����)���m�	��(y�r���_dJ��1�W��P9�k��9V�v����j�G�Ҟ�������'�o����-�֮�vAՃ��΄f�f�^Yc8Ju�"�c�G��%�
��>~��X�
i�O�*�i\�<�&.!b�#�<}�!1�@��-�|�L����9���u����>
X:Zԁo3L�Z�����D�^��d_�l�����~@��S�rqcӦ���b��b����K6�y}z����o�OM�������8�����Br�U	�����q�n+�P9�/ʆ2����[R�4�����ϻ?����jk5��K����+n0�ͧ�	ڠM��|@4�=g1�v��d�|[T�����;�f��oa":�Z��$�`��ι �6Cڑ����X�k�";�x��I,���i�8R��)]���T�E8�o<h�z&���x�&��'ΐ������ײ��[���2�+��m�2�ۛ���R�Ac#����G�6R�O�M�%�������z!�5�$3Q(���Z�c�����{����e�&��\&�H���@�zb_�n��^���H���<��]��(%Y�(���Ԋ|0*����S�0&ާ]�����C`9�aփx-~
A���=˓W3�����@�k7%Z��i�*M���`�R���:�k+L?���T�N�%��[z9u[�B�>�A;�%1�M��s���P���w؇���E�5�|U:%����>TT���my>{,�����t.����+�C��.	�p�*��֛w�����_�|��>�!o|bj�V%XF�fí5zxp�ia��A��Bf0`�v)8�����+��qn�D+=���նNQ��)��EQ��&T�p<��4+k�x��nM��L����<��6?
[1��h�$r-�="?� `#�L�A���@4T�/�
)痜m�_�k���YsD�V����AE�P���s����3vꘞy�����?��b+���:5�Ьԏ�� �%5M��6��1_�$�-�sm��rTg�,l9E��2�(}��?$N�m;��$ou�ǒ0!�26���w��N.X7[�9u<�%k�=���$(۝�`c2ki��4��3��3���a�+/�����/�~�t��~j碲d��#��6��S�N�g�>��H�Û,)��2�e��a�C�c�B��K�E3s�CV�PR�ݐ��mr�r`x��Z�	��P����;h����J�
�E:��y}<O�-�����X��l����� ����e��gs'yV�.o^���Fxg_c�2
�@0�O67�mQ�7�����~�6#�t����� _�껿�+��k�����P��bD�U�ȚĖ���|��f��4��Je�R�L?�S7�(�rP���q�fe&��=iX�F���K3����D�rp>vM
�\�eam4���X���r�K���+����<l=�`�@�>^����k�����5Xw�7o�#��K��
ՕDB�c���3�ն��X�-jz�Q<=c����4��}=�t�7F��3�ɲ�`�/����܏;�P9� N#zⶒ�u<����j/���xܙ�N@�_~�k��aR�*!�����Ғ�)��=�������X���y���o��ȸ���F�sF�N��;�,��������zʊ �$�Z�#8P�L�����II#�䶸C@�+�I� �U��vu86��y�f�~�2J���vy���Qٕ��%���o(J���jZR��ekx#�N�*�7��T+�	�	���Uav������:�L=�-t�G��n�R
ƨ(�ށ����0~�F`v=@�sL+�����c��zx�d=ǆ�z�Ri�L�y(��B?َ�c\C�ւٕ)tx<�O�aXNmXa�
ZL%r�s֔QPdW��쓏\ȸ��.oq;O�*��.q/T �guW����K���u��n��]ѻH�ke�i��P�ˋ�*Ƃ��*���V|��	���R�I>Q���R�w>��c�M������z����A�H��� ���ӾOks�1BCi��� �蟥/�B���9\6�N���ۄ�Ռ�*;|X?�~ߣ6�+�l��8�Ba�[�;H��� ���[ul�EE����[z7X�Sێ.,���(m�8<��^����l�˿����Gg����u��K�+џT�C���u�X��@�T{�V>D��V"�1%ڵ�c��l�a�?�$�,3��g�sRl�#�Z�ߣ�@�V�@�Q��]��l����Κu�|�Bx�敊�i�9��|�ѯ��; ��/C��x$�6,�KcҐ
6mdI��myWC
��;�H��@�PZթ[�;���7�1^2LA����P�&&��-�D�\j�ւ�N	��n����nO5�c�S�	�����Mj�?G!�<��Č׀���r~� �����<�*v���D� *�(��@��\���;��.=��&���ղ?Wñ<�$�?��
v������x��tP�d��N�B��W;��㲥�������kL��.�j	�Γ�YX[��q��l�g���Q��7ĭ#�Zd`kȋ�[��h���a�~2�g@��q���w�W#����R{ܔ�ٌ-@Xk����<ȷE��֖�7r��r��$I���ϳQj䝉�$ޜ�2,��t�,C�Ce3�0[ժ?. �11��$����lt�u�+q���:�>u�o�ګ"|��䌜#t����B&s5��_��_�m�L���S�����8��I�z�5��p��dR������D ���Q�K���[�
�-���x%�zc�Z�ux����axxH�JW���^���@W�W��W�F�y�4�^YXR4����n�M�K���a׍O��M��-q��M�M�R\�)���)����lIUm<�"��\�^���g�P��%0k�F���+��h����y��6=���D��tA�3V�#ZIT�qM37�᧟�_]+>�vh�L��!M�ME��u$s̢^�®��k���,���(&lK㎾�� �����/�y�Q���D��q�a�#��ؤ)20�˂�ӥ�Z�7�gqXL_+��4
�R��Ʒj�&z	�#�f����Y�����h؛�I���2�Gj�t�[�S�	�&K3�;��wR��I�G��i���Ka��~O�W�F���j�*�H:��1�t(��]O���ɪ|1Ei[k�~_�R�B�U�W��-���L��)���E*�$�͗��1Yx�V�$+�G/ ��,d��g��'�/���Cܨ3Ůn_(\�J���0Ĥ}�.��f*�'�\���3wl�4�����\!Z����{@是�(C��X���on��pR���Ǝ�c�����g����� �rf�o�EGx0��\�� !�������]��UR�±�u(���>�p4��9�ib��"��޻����_�{��ޙq�E1�M���^$�n3�r�b�@�6�����&q�u��0�PI���7�?��n���H#P�.SH :�5g���C	>j�=S�+�B����7���.*t�ş��rX4M;��Ρ�S�10T�jkk�j�]�I���
r/�R��[:�?�M���^7�j��D�{c�I�p1\EKÆP�i���6+OmW`pͤc�rd��Q�<�Z�eyB������\M	ң@ 
K�]�qO+�)�:W�]W�r��0��d��k�S�ʻr�$����������[��9�2�T��nWJ�3��JŜl���@���"�����T6�)��q�4����|�tC�Uyl��tm�b��9;�9 ���j� w����q��YW{M��ۅ%� ���u���D;�	;�DM$�����O�˒�r�"޲ή����3 �.��4�([�]E�"�����e0�����w�D���(B:e����f�R��_\�ܩ��T��a=-��Xb*ʥ��||�KS��_7g 7;�~g��h,�b&�' ���<��ܝΆ�v�4$R�Ү9�͚��ob)%
�>���2�����d�r&��������M�p�^��v��јjHw�-���������I��R;�����[��>󠲽_�<,����fR����P���ފ'RT�m.�j3W��Mّ�_��Am�d*c$�.(���(}��1������!s��$�{�1��aW\�H{en1�7
t̘5�^	�Y�;{����Ls�����Z�x���n�N����0,��ц¨vJK9Ͽ�G��i�j��aZ��"��D{I�م�Xf6�ѹ	�VM��+,ܯl��ᅟ�KF���>��Ic�Y�[��@�Ȕ�@8=�X��p��q$Phti� ������m��Z���!),6X���[�o�"��	b�~hߗ���߯��d��g��l�-������j�a�pBQۜ5�4�����n�W����ȝy�TX��&����i܁�TS�y<9<Il}dpT���(@�,�&��3��/]����Fl�.8���Γ�¼l@��xmt`����W�<Be03�̓���zݛ��<Q1)&��ȪJ�j�&)� >���|v���Ƕ����v�T��
�QY*桽)Iw:�ʽ�٦P�ߥ��֦�Q��td�_���*���1��KW|�\숼Ei��Iuٖ0�]�I�$��n�������Q�@{�$���-��[�k�����-lP��wq����ky�Lu��×�"H�������n����?׭�>�B̥g�l1"�n�9E�jn�����ה(=D6�O��CL#���9%A5�4)2@X��@ٔ�rf��?W1��=� �2W��Q6�S����r��ۡ��������h�-�U�;(h0�Jҷ��M��˞c��診mk(�hk
q:]���b��,�ZNA�5dh~�I6pCVPw�,U�0,O.�fpj�"�O����u{z�ĝl��ss&�	=&_;���Cd�{�t��Q�b"f��m:M ��}�,5�"�x�H�J�'�"�$r��=��B�C.�O�C`V�X�nr	��U��dvk�xr:�ˇ'���$�[0	v�-#���U���kЄš킁Ph���'���$򾌢�ī��pF�W�Ք`%b�Sg��):��(�	F�j�<ؕ��� �ET�H5y�� r7��a��kq�S���z �_W��]L$�z�wU�z�Pڛ]�ru�3�TK6Ĳp���KFV�UfU=��pV��HPn�����%O���N�U@D���eң&++"�q��7s�EsA6��~u��3*Z4r}����ڟ�&���.g+ѥ���;?��~��Г���$�q�l2�}���%�d�Z�ZL�]�C.ۖb���q��z«���_	��ʷp3�u���e�c���u���i����(�'΁&�����/Sv/MLB���l��IW&R�,O7O�Īu(���w�撶_㎄��UX>�"��C������;p�I���J��X$�6�Ϭ��LY�����ĨP��e��8F<���?���щ�-��HR���O>/.��M7#(���TG��Օ�[ptv�r�����KR��J��4��ҕU�_���󽄻 e�ٔ
��T&�>Բ�I1�����g��C�C�c�V�q_�vB�eo���/��pAR}
[i��}	�9�!L�s�+�r��ol��տ�b�H̨�Hy;!å�;'Pk]��hB^q�"�{b�*&���~�#Ϯ�����i!�ckt���{ܤ���~X�y��r>�9dq�7r+fw�����W�����<�5�t��J��v���UɩPߎ�����c�#���"���l���
_�Xp���@0�.�˱_�G����TCա鸡|��F"���R!�<9�o��7�ZH3�����1.���v��5T�/2}���K���;�X4��L��7t�t�z3��C���}���� e�x�o��}n��/�
E��ew��|���!*�����v���^	/�x7�eI��}q��Z�0m�y�����[r�F��"�����_����Ԗ
�X.��d��n��5�!#>�͵��OZ��j�&V��sǝ�$��ܡ�cA�1��W۰S)�1�M\&�F=Y~P�3g�1�� "�]�޺W��c+~�[>au�M�j�T˼���A?Ϗ���ۗ:�ˍ�|��p�`j?��Go�h�����*W�v��KB�Ґ��<��Y��;������AX%��4�5��l@Ja�m�	-�����V��d���fAy��H��v��x��>�bOt�	�)ug����Z�2ҥ+����	��U`�w�^bE,�Mb�����U;���Y5��"r�[(��L�	���
w~Ⱦ�IS��PBx���B�|��1w[P.:;�7��[!�H{�>��a&w@�cm�[:R�:�*7+��o�ۺ�_7�����?lFw��G����Ӳ�>��xv2���������B���}��W�(Ddd��Ms����c����_#4!�s��X}nİ�.A�Lo�l�\)*�*���:� �3=��6�Ȩ 1,���S3�^4���y���C��[�D�"��y���du�0�92�	�V�tD�I��q�_�v��Ԛ:���;��D-�RU���+N>5K��/D�#-3X�J�S��9�x9�w��2���:����L��ga�Cj�A�_��я�C����@dA��7�|�j���
$����awו�<�.Ĵ�[c0Q��r�����OwƸ����\ͪ �S�%^psB�\�(��9�*�<p���oe��qB�
��t�����I����<��mF��W�9��]c���9�A �
��/L	_��C�Z���<~�T`E_�9���pO�ų��F��L:e���9<�m�J���/ON�d��i݉�6�~�~�#
�gxi/��G��K�CѢ��W��뽡�0�V�@\��h�)��w�T؜l��΃ ��:�-�w�̗s�l�_��S�t���d^w�����K�J��*�^x�*��6��R<�)��k���(��J��k�^��	�4�C<��J�J/�xup"�,F.C�J�������Ȉd��s���I�O���ִO��'����>�<9�T���ϵ�uG ?�Q���6 ү鉚D8�i�G�dbp�Y������W�MY�'#w�l�^��Oi�������eo��z-/�sS�}l����;}Y�y��Wң�J���&E����������kFӪ�V@'J�cH-G��fb�m.���u�ʆ��ur|����r����+�J�(.��Mv�j�6�,4Q���X�>�5/@ a�`?I���R���сq^4���_�i&o��&pA��1FSX��K�duڝTͩ�׽��g���`F��a8C���t��Pu��=��F��'�~.2��k]���²�J~�G�4�������ğį���7=�I�ً<�F8,�=�����
����$_]��Y@� �Ե�oҒ�E�j#$s�_��V+ϝd������j��O�����2���nR$9�����jW����\�?N�=}uPy��-Ǔ�x~�b7XBh���_�?���a4���?P�����i���HB�Ўy�َ��nèr�n�%��s�%7�;�R����ƈ��6*�5��ZW�ׁ����dpp"��)�49��!��+#b�Ŝ�.��'}�/�|��{���ӓ�˺b�̲aj.=:�lu}_nCU/�UTgQ"�B��2�:��fo:@�T�z+gH>��3t�*��=�	J!�0���~Di��A��Z��2E���:��zp�F1R�b|���λ��<�Ϝ$��>>B�="�O�Lk���Er<�( O�9puc��C�׎�ኊ�§C�b`�cϧ�Y����d��<�"�ex��'>]m�gYy=�gY�1�&ЋԍWh|R lpbF?uT
0���f�|�iP�QFn,�G�'�mib��_�ot���T���i�$O�ͅK�tPu����H�q�"+ṀF5�\��yz]R��H���-bw#��Fۄ�J��t����s5(<�b�!3��P�뚀�'��Ge<��!�>�"�Qq"��P��,�+aƝ:_��Yho���L�f�S>���(7�L>�!��X��x�Z�]V�W�:�kk;n��f�؞d`[�ӳ4^`j�P#V���'$4�����j/[��$U��4�]��=�ѳ�'�0,�*5�_��|�hdM��(���z�5O8�P�	b�!V�S�L�X�+�;/��l%b�H�9/�
��ׇFd�>װ�H����w:�����ro�Qӹ���j�Z��i�ҷ����A�eD&���\��MX�/T��9�j�D
�L�ja�������~r+$j-��[�Z����B#��m
"��̼�]�'�Z��U|��X�����%�r�����3N�{1r�h�~�~���[�c�'=�u]>�� |3ԨDN���s�y�����lbA�c���=^�W�9P�g��)>|�",(o1�,n���Dh�S�i��$������"�0�M��*\-HE���?P)�{*���<K�%��b���4<N�`�1�/H��b���m/����C�c��1���Tv��iK�s�JT4LH.򮏪v�&p,���J�bba��^�g�d��&q.Y#AO��.�Qw��)�� a�ߊjh�w6g���@����!�,�������bR�n�S�Q��)�G�u�+���a�YY���\�ʆa��̚�!����Ae+\]��O$����=8.���~E���72Ǡ/�C�32!:�oy�d��+�k"&L- J�
Yv��$E�����-��F��(�"?�7��p�~�!����˽.���o�]���:�<�o�
�ם`�%�t�(�%��9H�l'��l���Q�ْ�5ͷ�B�k�ҥ����x���·��!
��cl5�A��[\T��[DP7��U���B�͸P.��"ieV�si�6+�.�BSx���������~R~�x���5#/��=,6E�=N %��&'ׯ����YiD�;�c'Q�1	��8�o�1c��3���В�JRa��ƢQ���F�!���IQt0��]��:Z��ʇ�[=��Δ%h�w�}�Od/�8���a0�sʨg?�sHy3�5o*��0��w�Lb��~�V��7�İ[2��O%W�n���"�jA�Y=��\���/����Ms_)B/��=fq��ϖ�v���Μ�}�=*!�l�E��Q=~�0DIi�TNi�L�xm�I��-���1��+kM�1Sݵ���>:�p���I4sF ���J2FJa�<�e���t�����߀��S���9�C������[��|@B���ҡ>���f����ɫ_Ry�������ۦ%X=}��{��'~7��'xV�7�g�_F'��ܫ�#���.'Cz ��Gy�AE:���tٸ����A-����?	_�ϯ��?/}�8U=���U��\Lr;���{�D�-�e`���3���Wj$8.�NRo��U[DΖXbYR�s*�=����N�"�X��*�ۻ��{�@��W>�ÑZk�9��P�˅�~�� [�-Q�N�QK` {%Uv��ڢ��X��O�[0��a���t�jބ��[T0-��Q��o5�Gܭ*6`HD�C����
7� �����aǚ��������q%���RmmA羹Z:b�\3����< ��~΅��4s��X�ybQc��:�-����6(c��S֖驲	:ǵmr{=ݏ�b�L��5�D��?�v
�eԊ�� A<j�xm�d)Β�����`&�ph�p��N�gRj{�VL��K�ef�u�{�c���̌�n�h�f|R����w)���@���u���)ߵgf���7���p�2*)��N��z��L��w�q3!��Z�_�9�3N8�ެ�
�1����ʷ��/�Gg:����N��B��.m<K�ͱ��n%T&�K����Ȱ'���{���ۼ����*��N8�E�.w��<���!'���X�_�F�|%_l��d�8�z�M0�����V���>HdB��
�����p)�O��L�Gn�[�i��uӥ�R��p#Y2m<���r��F�+Z�G�om f[:���\��뎒�|ӳ��!���d���U����](7�67G/3��#ѶxM�����E+��|�K"��w��B�\:y,A>��K[�Yk lf��� �T��PbF�d3��?�W�_P|U���)$ѝD"��R�H
6�Uo���ː3E����h �{�j��g�3`M�6�ڮ��{x��;r,ܭwۉ��P�5V]��)��7�j�5'@������Ek�rG�5��>(>v6�2�iKHS��F������@^>6�{d��
�@R�(C��~�� bˮ�,�H�Q�Yd"��J��O��ɉ��^�C�EE��4��g5���1��/�����
k�L�|�I�59�3y_
~��ts�Xث���O�.r�Ę�?J�Q��S%����#�����/�w���j���3��������j*H|$����Y�G\K?񞄸��A�>��Ki�k��
e�B^n�{��o��]j�>rd4e��i��lKN����LJ/�A5�p�֎j^�sp�V)�m�١�M��Q����鏒��9��G=B���#.��tAն�F��?Z����8��D�
����)�B>���|v�s#�hD(��eV��g���Ŝzgڙ�$򚗱E�P����;,<&�[�,������o͵t��!��j����a!Y-�aG�t� 1;g&\�q�����$����n�K��iY#����3���f9�⨍�[NK��Y���f�`Nv�a�{ �4�)G2��a�V�	EfІ��o՗���E�}?��>�k��0T�f9��������݈M����;-'�-�1py|E߳��D�S���2Φq2M���:�p�uR}@�>����H.d�E
��d�g�_R[�&V�ꄇl���v�i��]�m �z� ~p�H;a��WoKA9ᬙ~�ZyN�h�P!��:뱃�Ȓte�Ӌ�p�K����\0���4�J�Q�a��p[z}���CƮ'��|,���E	�j\�ȷ�؋0s��� X�)�sL��4�)����t�O�t0������)��Tf28�nMk��w�׽��J�.��q�A�KKWk[�1[�!u��۹Pc\ު���Zٛ�V�f\sގ5r��l��>��0���H�o�������N-Ǣ�M���G��L�Á�R+I���O�j��G�]��lò�P@ ��r ���W"��V�1��\cQ�؆�,ܼ�!$��W{Bg�?����q�, ��DL�����rtuϟ�g�U�B��="%�3�l�:K��{�?���X�L�5�Ե�������[��ǻ]���ӈ%��oT��0�b������"�A(Ļ�?3��a�~Y�����i��w�6�/�� �̄	�d���Jgz
�\�P�\�f��(�:{
%���yz�VH��o.?1�F�Gx0�*Nbǻ��{x(�ky�d���-�j��eV/���
���7$��������(:����s��l��8��[��#�:un_���`��-�tohI�V��ӓ��ǥm��rG.2-��!���Y��C,7G�.9���#�+�M};��G��2�I��0׆(f��[vf�)F9� ��I�ۼ����s2�����:�~�J�S\�tۺ�����QA[ԕ����D���guc�x�����'�}$�*,��m�I.]��Iv}`�,6RXve}�W���Hqz~�F���Y/s~"���T��0_^�cCF����˖�6A�_7+�o�V��e�5E/s��I���g�T1�����Z³1Ȱw�L������$`  �ڭl\��C��'�d�v���j���χE��n�f��"��8���u���@I{K���|<�t�Z�����9�s�5��3��~�Y%V�CW�� �4&#��^G;b/���XOAl�� ����F4Bҫ�\�6ї���n�{;�=�B1&FTlZ	ph|ɿ2�Ň-�S	o�5n�
 �G>*�+�M�������+��G��ɉ��g�q䞄�Ј8H�eX�y���R�\]����R���߂涝u�U���P�]�BbJ�Q����o���Nܓ���s3���? k7`!k��8�6jw6�D5�%rMr��,�^�>�扈����&l��*���"H,����Ze��7��p�7'y]/@p��'J�"���g'��f�-�[������sB��-�7O���ઃ����KF��0���強�_���b�o�n���}�e��x�H��V��``G?��}Ϗ��KB�C��q`��Y�eV��q�v3ש����@_O5��*�� �j�xC�Q�e�ȱ�.��+���d���']��kf�@����B���TZ�j1x�k	ca�d���2Z٧c��'��,V��~ϼ�� o�y��NI�5��Pmyg$;���w7�A�R% sx�wc�TƏz3����F��s&�H5��B���!*�>�&��o��tM�*���E���AOj�r֏['��K�0ZZFoA8UR��}��)��_�,5?�T�.(�Q����̦T��sbj�4k�q����OBq�t6-n1�yU �w9�h@hȲ� 7?�g�M�]ky:%�.�aU�=�v�����d���<&���� Y����NG�k�?`f������O���?Fq0[+��F'y=w�\���0�[��J`+����,Ĺ�	ť�|)�-���,lX3�G7����V7��^���;�yۋ�M��^ZN�f��6Bt�p<2Z���:DO;	8�4f��h�b�&�8���A�a�R|��IM�����dOž�!��$n�_�`<�3�\���+T�][{��w���}4��
Uw���>2�1�}�H�S{+1�Z����X�۲U(��@��؍���Rym����`� ��;�!iJs����`q*�n�`;oUX}�鴯��x3�7l~��g�l�b�Ͷ���\uT����>Xןs#�	�u��u��$�9?�sv�'�����6�>��%K�{�=�=�尓p<+˝~$s"sNs[��