
module NIOS_RFS2 (
	clk_clk,
	reset_reset_n,
	led_nios_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[9:0]	led_nios_export;
endmodule
