��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%����씤���uG��uzCOkK�A�F�l<�3$~�>7��D�!ު���ő��3 He]�J��l�ߡ, �
������q����3q�
�5{�.똴�l�=)����-E����k���IՋ>����|�Q�;
u>�`1D|�F���l������m��ge�z'U�Xb��u�Y�z�3Z��˧
G�e.�I����gI�a�XC5b����<�-'A>敳�f�����)bT;�h��頣��tEUޜeSŞ�v���Tb�-��J�$S�� ���\����F�8m�el[��W�2�M�,�s�kSc!��U6��L�ROӴ���CX!�~���SJ��"�pG�����N"{&*m,�A�/bӏk�0�xM\��[N2���Z�kazzH0����|�i��	�R�&������v�Y�u��2_O�'��p!C���+��a�j*�j{��m�-�S��c���gt�8f���t%��/�S��M���[w���I�4��a߉h�[��'F����w�������������SIi[��u��X�phB��X#�TI��C�F�R|�WvXu��<�4R��§�܄��Sb�nA�4�Sk������#�ɟ`���-�I%�ȟ�LDO]��c�s��	�z I�ޅ��"�6c��\w���;��`��r	��9��q�{Z�?��8����z&
�&HK7c�jO��)_�L*��݊^t��Y�h�6Y�b��m���h���oh�N@�Wں�(ot��b�6n����ZR�ێ���������C�0M�����Ą�� ���bc~��0�{��/ww)��9��SL�∶q)�'e��;e�X�MAUɟg�ԃ�e�$�e�ϖ����^���W�&{�����(��7���U�4U�ǚ��E@Yg��W
x���Eiu\��{VD�v� ���%>�A�i��+���둊69�<afjR��Byh�ߵ�wV}Q�20@6�7}s�	.l_�R�gy��l��B�{��p>�WvnY|��ɕk&P��U���'��������@�R%G�M���&�����DSeU��<�w���l�m����V��.X~�����=�6�lYc��bvP��0�獧O3\j�R�?d� �T9fX��?�o}�8�����	������3'--_��ĵr
��z7�csB&�����5y[2�������J?��#m��D"P�Qӳ7�3Pbb�<�s�%�a{f�h��v�7Yb���.�P`|�=.�|S���5�ڼe7�c�|�u��H���>$����!��P�P����|k����2��,H挺��D���hb:z���.���_��T ��v�[y���"��Л�ZD����J�`�y�JD�{k&�d�7��/�#k��ְ��'(#O���<��'CJ9�¾@�s�o�ё]��r��_�q��$>0�}���������{Z=�������*캗
���5����f��򗒟j
t��ng�z���D)��j-������x��|nw�0�Ӫڪd�](�	.�"Q��EB��v�?����B�ἐ	�O9G<W�d_�R组9�B�\ �vr��fC�_�vW����e3��Ҍ������(�83sٺ�f'�eG��d�����W�-��eC�T\�rF+���<!��~̕�;�$#�71� XfM�wV�h�v{ֿ���3��+Hb�x�.�+��%(ψ)Y��\�+�ބO���g�kD�iH�t�Յ.�թ��z�X/ d����� D������Ea��#��q���vF@A�������U��aP43Q|F��Q$2ԩ��J/��ԉ��J4�+�e��2�&����`-ց��/�]�{�r������ٌ�������eD�'�����q��8w
^�8,������J��m�KO"X�)n���|��ICf��`���_��߷���&��y����;BqtǟOAZ1��.�fU�ól�+�k�`R��z�#������8�T�?��*R���g,��Y��.�ϕ��	X�Yr؄�V[�9�Q�I�8a$X�!�.�J�t��Z�)��{�tw��7e�!�ľ�'\i
�E3R&���$䀆zG.H��'����G��7W�@~�۱��ē�៬l%������W����pT��xR�~�� ��'a~B?L��L�����#s%�mY^Jq����UG�_��X�X��T=�m]&��ޞO	�a4c��Ģ?��*�T�x�M������%AO��߽^SI�#x�\0�z����ߢ�x�?�͞�[����&��'$(|���f�U�e��;��HQ6�ϰ��!��i���2�C��)Gdۋ���mU�.�T4}K���@_4Nnt2���������-kd�heDOq�ᨭIY��s�H.���x~�k�u;��lI-�0��j��&���nq�_���J�;���l�9s_�����fY�rUK*��b��7�0��U��o�S���,�0�8-������g��ۘ3O6V^qn�Qu`'�l��I=�]�J��_�Ʌ*��12�{.�C��bW�ڰi����jR�*��Q��kXU	:Y�o��B�lp��GA���YI��Č�v��P�OZm1h,r�8�o��,�+>5y�����\��'Ժ٢��$.�)����� l؅���.�Z=P_DБT^�V;������o�,���'�v%Z�L{k?Cs�
�dn	��W.�f�>D����F��b��'I4�����S����B���gg���/�����k��+1y˞D�>�*�_ݒϻ��7=��-�xq����*��Z DB�/��&�*�лI%�0m;�d��yM�"��9�������5;>.1$�c��4��Q�c��o��f>���;�����Φ.�@��W�8�V��V�(:uB���r��w5���%N�(����7�s�G�9~.�	G�t�^,� ��3_a4zC6v�@� �؝by-.v)��i\ ����B��q��pUzC">�΢�	�������t$;}x4%|���~�\��^I����r�>���ʊ�<ن�#�H[l��f���\Vk�<���W9 �=ueX^:�������QZֱӛO�p5`�Ax��4����c���n@&@1|�2�'J�=%��oqz�M�xB|�d��0���N`�#�y{�ޟ�h���é��a�NX �����.*_�S��*�E�ub������K�4K��,,����,h��=�)�<��)�n �����"��+(a�Q���a�2@����GTW���Blb��b�J}j^��J;e��^�2ˣ���YI���Q� sN2���shb��Lɇ�4��m���s�՟n"�LЍ�I�蠩! ����5��Z�f��f �2��;��� EN����ڐ�Z�Ѱ-k�HV�ň`揲l���f�_?jQ�|�:6��J!��AZg'w�w��NC풾D�s�0��ܬ����G�,��ږ���Jm�~���@Ʒo�$�nħ��5%�מ�OjuQ޹���m�»]�y���>�4p��*GO�r��D��XUY̠�;�U�a�����Iɛ�R��O�Yz=y@λ�8��:c$tr^���~$�k�������cM%i=Pʷ��X?A6�UR�r[%�	&�H��i��R���Y'Xqv��������G�����bog�9�`D���˫;N|I����תƿ2�5ؔ���>n�3G�p� �㲣4 ���n�z�ϭo���
�A�rz$�'���q\���I2�f�N�X�0&T�U��\U[����	�B�������Ȑ� W ��[��
�(�����ֵˈr$IK�	U��;�?+t�j!�\�}�\�"=̑?����d[��5���峮�����/��k	�OB���璵^Yr�Z���W2c�K��\Q�Vz���AXT#Z^��,.\</Cj��	����e�]݌Aկ�X�s��c}
��8��Z�+;mw�7$: (U�^ַ�ڶi�w�J�u���fqG,��q�ޗ���_~��zY��y����ɒ��n���X���:������؍���g������Zr-�z/���4�@%aO�P^`��v:��A�C��Q��!a�pq�.��4VNn��<<{(����F�r}7Zh��K�*	%h5q�ڍ�(�Y���Z���\�E�rBP�ks�R���' )�8g�����ms�%��|$e,�ɵ-��m��#t�;���38�u!�.��b]P���ԥS*�y���:{������M
B{����{?'���nGx���&�Y�@��.�	]�]z�n�(܈\;ʯo�9`�N��ҌbN�N��΀"Zf�B��a���G �'wZ�̉v{�v;*��Io`�ߠ�BD��C��Q\_gn8ՠ�G�����طN���m_����<-z��V�rC�8]��(������	mh��Vvd�I�[��R^�s��g���B�(�tIP���f�И���7VM���Z���:�ѽ�56�U��mU�s�V�	}��=�:k�o��B�i��3
��،6(`�,#M����	��|��gۣxl@u��u�8��gÒs�˝�����
�7�>4"������ s� E������i;�sg�d��?q����،H�Q��<;��6��?���?e&Wm�J�iR��(�hz�|"�M�q���I���>v�3h��'��e䁔�U��MA�ջ���Tu5�}#��,� Q�����w���N���X6��!��R�A�>�ŬN�
��Da/��d��z�D+��l���GE��ɣdU\�;b�	��w���M�E%]ņ�������]ϡ&��#�^�".6�A-1c@D1�h���3���uxM!D�h��|nm`������I�lY6�dIj^��ZU���5^EUW��!�u�+����+1C��[u��>$��ZۀIk�C��P��xX�M�II�i����(�`���]S3K9+����j��cs4�Ҫ-��[}������6C��E��e�x{�].]t62��7��meMԒj�)Vh媦�����{d��wx���A�c㣸���pvF��� p�'q�ɯ�-M�k��Q�:�o�!H��T�a�:%�5u}�%�B��s�9؏�R	h��(	e�y��
�K����.�����d��$�o��E��6w�^�b��^l��d|�KP?H��W_̎s�$�0	m�e���n�1��e��$DQ��蟞-���E�N�J��ŝ�1Ύ�m�� _5��|�q�����풴D;z�q@V�^}Q��O�-����'���ˌ�a����a����X��u !��hp�S���l���V�3K����u��8݊E@���AwP�
�57Gұ��/˂q*�r��}�I'�����EP9�؁�T۫xW|�H�@G���09��yZiG�X�إ>T H��!vף�g�wo�k��&Xaz��a���-Č� S8��R��LDI��jةٌ���ȍ�Au U��A/�I:���������e�yȦ��
@,�����aC)mRX�&%'��H=T�N!��B� ���R:b�e����������V4��FOl,M��銪�$�ɼ�ݵ'��̼?��̴?o�|���粗1�:�ߛ�����D�٨�Y*��wS�}�;���<�\r�Oa]���%+⍫�ʴ�?GT|�J�s�kF&��ZZ�/sU��5��$�^�L:��l|�!�@`�"W_*�Y_�^����M$����T�o5�.����l�{QI�mf6�g�~�Ȱ�nZS�x���ü�?�_;�Z��kx\�@0��E���?���@H&�$�-�^wG�#�,��l�*�&C���6@�e2lH���������g��9<j�ڠ�E�X�N1.��ZdT.��d�>�H	4�ā)�0�����Us��g�G���i�񪀖hDx�
:Avt����D�G
�����14r�xi�F-,��sw1�ne7�n{aEs&�H�*��(�!��R߾��(�.��`9�Mv
���ǀűfK�b`
���ƶo�a��p^"$>�9,�;�'l~��#g�
�m��5��������=�O,�����Ќ��YP��T�k����	����-ݎg-!
�]�6�x:��}��$v@�rs�F�zdH��[�^���������3윥ͽk=#ꃧP���F,.������٦3���C}��������FIY���A�A�O�o�
Rxky#�P���a�T�՟��T�M
�	ǰ�D�LE��@7��0h^}Ѧ�0�Mm2��5�G������QS�=���_�p�*Bw}�0l :�H�Α�����º����4�)��A\+z�;���v��D>�����8��������`]�]kE�j����p�*����B'��!Qd�D�Owc���s�e6g� wR"�[�e�b�ʍ8�Vx`�I�6I)��~�ř|��eo��:����{�݌4'V<GRD��n�U�D$=�Sp�*�����||��c����̯2�Zk��}� �f�]��4�hZp�qeB�K�x��+ ���x�Ei���d���;3M�d������k�'��E��>{^�)EQ�邓�Z4�.��l���-Z�Pz|<��뤚ɹ�%���:ע�&�}Bh�
Ah�@�	A@�3�w� &�W[��K�Ƹ;I�a�pKUw��V����7��{��ET?\�a�G�����"P��X��h��D��c6�%p�AESTZ��I�>vLf���w�_��丌j��ٹ�?���֠I�ҳ��>��F�Gv��[�t��
��<��g�i�Io4�G�:�:	�o�w!�I+��P2]ĵ0�D�ų�q�\��6��.3�T*]����QT�a���S%X�A�,lAf������Ue���v����(~�+G>AX$�t��~�\୥���P�������:��5Ϲ�YG��@�K�c����D ��+~��f~Bp�&�������{�c��qƵoyW�(_�I�g8�7.�l����+�uG�!>j����&v5�T�JշyZ��\j�J	��g �xj��L[��E�@�y���$ȿmK�_1ߪyf��l&D�����Ɇ7FV�Ȗsr�#U�
�մ!���_2R�Xc@q���Ջ����qEjB�d���9� �`/�P�t��/�6ͣuhF�]M���{�����}�
Q��Q�d&�����e�c��Oi����
Ub�u� �5��I�kàx������G3�m�Ğ�����ؿ�v�{��n&�4�6���n�g���	u+��3��	����'b���ЮZ�~2��r��	��к��;I0��"�}�ײ�+0����/� �[b��'�op�|�ny�t��9M�������qo�ˑ2�'Iq�fS�}?m*�Ž1��%[v�R3bo���q�)�U:����U]ey�	>&ɵ�;�W������(#��
V�qOd��P%E�=���儳�ysIj���G�)��P�?��Lb���	S�]n����%�Q]�|�������\꥛��f`Y�᜞�KG���d���W���P��joeE��m�W_�gM�U�΃>@:���W-w8n*,,�7�������~�~ ���I�^,6�pZx��_!�Z
��w��4�aP�us�>�z`�����m�nl��E቞L�������S輏Ѽخ-y�&��p�`��7�cu��SwC�-���cU���(����nn�7��?�`c	y�6��Mkx�%Ih���\	��q�?��zTU\�H���;�r��{��"kr�V�i����Wa�uR��qTo��ݑ�vI�?���AY5�LJP4���ы���Oz�E����8�1읲�Y�R���wT�}��s�=��V�R��)ػ�B\����z�q=�f��<��0�$���p�V4��8�r$[�.������)�@Xѻ̿���Q��Ic�����r���?-O(;���8�x�E�uz��eُ!���r�oqP��,U*�_�r�4��C0��E�gT&��iQ#u�ż��At�ǻ��`6~�7#p�3�G���|��{�~\��QV���^}��3��?��~��'�W�̕RNC	��X�7�4�OG��εtV��J��/rleKK
�b��Gh���?����7K�#��H�^ݡ�x�ՐI�����!��K�7�|Ϗ��ə58%p,��)�51�
�ֿV�d�9re���-��ݺ��8�ۙv"\H?&�{n�6�,M!ogL���ňL��ũ��Ss0>҆uk5��i�&�M���~�o��{�ZqJ��hT9F�Q2-ipt �f�����&-)Aޑn�̞q]��-dAz��V&�R�O4���x�w�c;��7�x8_=k��y�)<'�C��VN^�Q��}��0Ol�ueV��ri��<gfUJ<�%ev�Y�?��@ϒ�gQ���㷲	{k���φ�#�S���Gy�!7�����a�O:�'��z�-�����1p]i�b�8ǉ���t�ɹB�CFhhL�Y��ʉp�\� ���y/@�Fq9�ةdn�b�b��,�»s���KL�CbGk{�l���
��K]P�&�V��y4v�q�XjbVP�D'��rC	5�)�|���lR�~�j�2�i���4<4=�pp7lrw0�Ģ!ܶ�i	fA�+��&xq@�<�f����v�����t<rR���z<%Sy��(o��!W�j��Ṋ}��4f��e�������1e�;Nx�@��}�u��KD��x���
�BJ�X�Į�R`����R�4��x`X��<5a���l�]���|{D��v��o�(hA����?jkFiZ��\�6Q:ju��/س���C�7�qT����TKk�n0#t@r�{��<�~f��AI�	�I��y�>���M�$�iP]�R�3jʂdL�n��+ѣ+FO���p)k\k@+�@��к���ʄ��<��XSAEO��v�Ռŉ~o��4���+�[��
u�&h)N
��s�o�j3p���C.!7 �[�v��#+�P}���T�:hL������+V9�����۲;�wy+�r/�ƀCaJ/�!@i�>�h���[.�O9�+�56Чg��R�$;ŉ(�å��ͭ�"�|@��mV\���t���,�����,�6��G��9�r���V2%������	�n�Ɗο�-����s��HR`�a���1��{���$��8 	�ƥ,�}�t����SFSOC���g�
�Bef��sI;>˕V����i�����x"e�)Eԧ�$���$;�1~�}|���,��r�(�V��eR_bSl�5m<���B�c1*���SF�lp��ًB���Q���^�^��c��_v����
ڼ�A��X�D/	H��f��W��I�z��q��+���}�14��:9�.���	����?�Q��BX_zz���%�d�E��zg:���L�pYg�Mͪ�������J�Ƥ6� 47J��٤�΃ə��!!5gdm������k���o-��ȧ� Ú����b�>�����qX��N\ a\�Kj+W�)wgE�!y�ӡn�Zml��5Ì8	��#���/]��E�<$����3<ݤA�M2lA�[rV �s��]o|�B��p�7������'~�x����zgD�&	e��h�Y�����ϭi�����&Y d�r�X
_C�M -j�߬��"��:���b��T�̢/G�b�k&4mb�+�#b�9A��D�޵��S ����Tn�d�G/��>c�D__/Q�wI9���*W�� ��Q���2�����t�V�2;^xPq����웠]�����E
�Զ�����ܡ�E=��?:��?������� �<�yi��rc�>�E�!�{�y6)ν�.��
(���Ss_c����L4Y�(	��0s�6>r����'����]&8�B�%g��b�_�w�,���$7|�����/�R#P�1����*rw��s�!2I��O+�;j��AGjF�(vD��z/#�x9�p+�	&�p�d�*|3i�Fף1��g/zZ5xy�GՒ����Fd�u8	�~�':�S'T��c_��?�01��]��}�~�x�?41$#+o�Y���`�oBZ��*���l�����⦾�a�@����i��?w�`ó�)A�e!{9�Gt�S�
�7���H�Ȧ�#O��f-%5�~�u��5��}� ���!j���6�������.�i��v���E8`�	s_�!x5h5
V_	;8`�� �":��_荿��AV����P�nO��/����<�bUw�?*H�rBb�n���m0^2k�E��k��Σed����o��"�%���s;)�s4n�`�:�#�>Y�Ku0��vJy"��v�����x��7rg��em��2�s���.QD!r� 7����2+zSY�(�) ض�[�&߲w%�g��2��<��G	y8�$�Q��� �W���CN_*�C�6+K�� ���s4$	@.�zLsS]/{0�P;ǚ;^�Y��������E�T�������c�+�;���C ơen����6���w^�eg�?)qn_�.s o�	ol�� �2�"��<B�F��@������)��Td�ҤY)ECt���M�gð�T��.���1���z:Ix���+2�س��c��-�Gp����'jN��hX�Je�'��ƕ�?z�Q~|�S6��}�.˯��e�d�ȡ+�0������Ki��=��F���Pxz������:0������q�yW/^���>j���jX�J�ϖ��Ic�K����֗�E����^��-6�qŋ�et���6�O�� �=�"]w�lU@�����)|dh�uڔ������U�!�=,gɉ����2��7 #V� �A+M�]�T��p��LbDIǾ�3=����f��8�}�4KQ{�����K��o�^.D;��k��<
��K���f�����0�vԔ?�����ka'��Ļ���Gzer�XI:�v���+��L�m�,��%���S�HL>��.(��z�(��&�C��|��z��տ�9v�,�Ѩ�:2Y��W���|�����|����b�����*�\�9���R!�Q	�D ,�N�(�@j�ې΋��ao;�?9�,ۂ��E�!����M�Hzs�����Z]o:I�޳:"-��ӃDu�A:�q5�h�n�4KVc~]�T����)�׀�|��*T(̤�^>~@ �W�a�]�z��a1�i*��[ ���^MW�ѵK���R�Y�%k�}u[�Z��(|��G{�(��TcO�^���y_-l�a��4U:�ke����\�=P��PPլ�kJ���k�;��@Y�by?��c����Yu���Ye���W�<9�F���G��2N�0YM���?͓~��]��;�u��c�x��O:8�=���MˤY�a�'o�M�9)ns�%*��(�4g8)}�#�
�<>�"_7��Tf>� ���4~[��ח1L��P�������r�̔<��Ji�.���*;t�dX�=~7c��U>���$�&O}�;��>}��7��h	7W�=4s�t g�����z.�Y����.�b^;�r$>�Sp�N"��<e��P�u9�)�o~��W�R��L(��=�
��N<��Rm�z�Ew�y���mp������T���+�￹[��>��_���:���%7�D.��_D���	0�/��}Ɓm�J�K�Sl�N㝂KLDm	�bޒ�J�},s���3(,O�Ά��_������L���n~�(�d����̎Lmny_��\im2Q$*	1��p��5:�/��4^j�:�#�i !'ƫ� �)�`q�}QX�սl��1�[���e�Ȳ�R�7�h��G�u�RM��(g3�P�����y�_ ��3��B�.P,����}�y�ʐ��A�9	]�D�j�UN�mIᎆ�\�ϊ4�v���7
�v=��T��,UA�H���3�(�Ž�d�6?k��h~�f4�w���.Cc�������8M�pK��Gϋ_к�d.�*�Oa�Gm�u�8#�9t�B>.k���d��c6t�'���F
���e!����Z�r �bK�f�K�ɍ�x�ᨰ�
����G�<eR�M��Z�7��U�,3g�,r����������t���^6������^i\�d.ʤ�ȭI�wm�ach)	IFP]�K?�*{��:��۽E	�=���E�_��f@6 k�a#�#R���
�k�u�g���:��b�ƏN��Nđ�-hT�@��,a�H'�d��I�G/^��yڙr���>t��&�<%��9x*�)�a�����x%�Qu������j7�td�+��qS��K�qV.��ݟ<�ނ� �[��W5���C��S['?��S�Uy|��d�k�9>ݝ��IS�6��ʓ����^�4�;��C�s�ȇ���l �q�ܵ4��͆&}��,�m#�v:d9J� !D�=��D��[�����Do2���d(~5�rW'&�˺�Ȍ��vp�!K�^ˆ��'��{/�)ݷ�2�:^�k�`���p�p��ilgb/yTy�<x?��*��G8\�,bJ+4��e�'�R�Xv|�H�j��/6���}#Aj��j}���(�Uy׷��*5$�5s`sA��^}T�q� p���>2�E��0�ٔO��2W����H�3�g��u���l�c��}_���ⵊ������h�F�k��p�!hRtúĴ�@�k;����╿�@�K��QM�GE��z��8JI���T��sd|���NB�P<
 ����Ny�ڸ��KŤ�@��R��=�t9V������3Z��~l?����O-�P���ӭ�&ƾ�gڬ�	�}2���0[��嬄yG��t�4�m0r���橇��p������:���
e������Ÿ��n8M���m;��v�+��� 6H��:�{�y�G$��x�A�[WV{�9VeD�x��2�[F�i���a�a���u���9�X�{�ޠNu�-=��k^�fԷ�j�@x�)�s��.��	��g%r�1��; ��2s�[��܋� ?�_#SNd��*W]��Z},.�7[Tb��		sb��)�$r�6Ù7c�)�:���l3�5˻z�q�vt?����yM5��3 �}��ȪM4���
"�k!՘�م�f�!������l@���q�i�e�6=T,�JI!"iN:���QJ���f���,Hr����[>.q�?���$s�c�2���|��P.�h5�
�a\�ǐ�^1Ek��;�����������n1_٭(�2����v���|�O���$����ڇ��n���}qb���9�Ɨ(Ra�Q���Q�o��t5��K6J[<��I7�R����K7HM_�����*�B�^�cEX'���k��`�H���%T{�,l��@*��T��E}z.ɇ�����q$$�`�	-h�$Y�%�1�&12��&4�C����R�G � >��OY�3�-��=��Q�ϙ��ϠK�Ȱ���YQJ>������ >20ڱ}�������@���W�����HS�)U�pJ��$�<���c�C�/����2%+���Iq�����J�b UA�[LA�,4N�uT�Z��+��A���e~��%V�)]��M�G���*`�Wn���Fzb(@s-��Pi�TPA��k�	��k2\99x	M&3�z�pi�����l�޵�U!�)��M�R�"{-�?����T�j<#����	���L�בw��u���?��$T�W$d6x.�曆���ZO%��TF�BE��e^4��#i���Zb���u�!>��S�t"�{�I��O���ݙ��~�����ez�� $w�c&q�����ϋ
x��d���	�{N~��Dw����^Fχ���&�CP�������P���[,#:��'�کJ�A�LU��fQ}��m贝 LSv#��giJc%9���p�
�-1G
"�@0Ug��n�@�u1YB�:�^NJ������{q������a�4x/T�|�~��ő�Ȉll[e�F�{�G����f��fO��X.�)��íJ
J<E��c����x矁����G\�G��>͒v稉�G��)s�ϴ�~��D�)���U�+m�g�+�a��A�'DW-:%qG#@�QR0�az��.���)�Wzm��I�t$�d���X���~h�`��?=T�t�^����T�(w�,��	8�X�f�J�δ���c�.@dj�X��37`s#���S�����!f(��I��r���I�����({��ϟ%�	�M��a�	
�pL��t_/�D̻�st�=�%�K�Ɠ�t��X�H���h�j��z�/��m@-/Tw\���{�0����7�6SCǕUQ��*��'7�谒?e��fܜ��q�5�6DylcH����Y��S}EO�z�Ӳ��>q��_l��@�C����\�%�u�.z��i���n�r�O�w�2�:�����!�iwE�^#yt��K�X"i�&�MZ-���zv�s>{��QN�? ,~t�1�*?	�+<�w��=/��F�B��9I�����+��N�Y���������Q�����a��H�X����O:5�2n�l���K�s0�P�g���A�S��E%���� �3i�t�M�9pu�q�L�,�2.H�E�T���ȇ��'�k�%V�)Tk��H�E����I�-"�}����dg[���SUgt $ �]���|�`�s�;�:�_f��Z�#����j(��͊g������=_̢�� �]�5";�6*,��m���w�|����b�m�nG��V2�������&���� ��gDu�j��O�j�T��+#��[��le;)��.�Z�Iք����="�pr�0�Z�?��[��,L��3�<�3��,1/n��}_�FUZ,^�LV�,Y�:X@R�7_�t>ؿ���L�	9�i@�qm� �U�B�����2r�MQ2�y2���Fd=T�Z-6c����. ެ����۾�a�_�}S����{~Bt�~#�n��q5��+i�;�"��*�$��*���n.z�A��c�~U.�M���Zr/^r���
�&�(3h��� �����yBֈ��(�j�aσ��P]
+e��[
����[�J������Y�ޭ�T'���hK�Le8����hF�\���x,�|8�0o��@f�D�q�n��]�G*���@�7<r�3�X 9�ʼ`lO�[���^qt���o=!0M$���%�>b^�ɼ�a~/��.̃��lyn�Ͻ�ZQy�%#��j�o�qC;��bɟ����e�^��V��ı�kd�Osw/�U������,I�1W�ٮ#ɺĤI�S69�>V~�w�P[/����_� �=��I:CA��XA \�f;ԟVO�@h|@�ګ��$��j+!gY��!�*��?V\�ŧ����-��S֗{@y��t-�a�-�=(	(�i�`�|�e5��35�B5�Z��38磜��p�Se* �iYLX�t���k���em�z���ĺ����R��b���o;�x�5�MC���b����,�!]6Jwb��'Ƌ�����;�?1ٜ<9�:�D�� ��A����K�d<o}+@-��T�|�tX���8�**ƞ?
�����u:����2��!&�E��~G�IFm�1��p4߲��7�C�Ն���ʚ_���6~�L�;�b[���#�V�� $Zṣ{�@�-Ʋ�{�@��8�iǱ
���ǡ㍵�A�`����1WF�V%���q�
Y`n�6����0-؀��<�<���ˑ��ab���0H�^��[�a2�P���i�E��8dvz�Ep��R�}��x32?տM�y�.mhӴ6�����ڴrA��j��ʜ�`�VR{x*K~I\
)�
�<��7t_��P共4�~���a:E�Dne�U�_� �,�%L�<�����7_˛n�l=r2��ƀF�{�sޥ�r��+��W�g�Ȋ$��l�#�_IM^6O�8q�Bxvńl��8��H���׸C0��=����G�#=�n0��4X�,Z/�_�Gנ�����"|
�:U���h^y�xo���d��R��I ��������<Xn����4�n�W�s�\1"֎l�7�/�����%�3ST��B��������������_}D�J����TM,.��[���!ӏ�p�X��D����'�?m3mT��:�qdK���g�!r2�eNH��;��� ���;�
�����^M����� ��K�Rw�';���B'/�jyc� ��2OC���	�Sc�,��-��8�5�C��Y �,�ȫg���g��S��>�&/�㬟�},��]�a�K�Z��g'#3lXP%}0u�r�u���u]�޶����%��PB�>I~ꋣ��+��m;�B�k�c�w섯x=rcD���f�3)�j:a
�k��Y:�о�)k���g�΂���W�������U��l��Q[kR����^)�R�0v����HY��Τleg ��52�1cY�M��:��4����śj�φ]qyµ�0c�0�m�y���CK�H�Ƙ�79G�:@�+1Jz_�����%�e>�>ٵ�F/۾�7g��C ��($@;���j( ��6�e�7�����g���p�M6>O�'��q�A
�q׻o+8e�4'���E/���=�A��!�To�먺�L�X+[T������H���{��;��}�"l�݌�A"�2 8�8��c��	@#P���xj��9z>���U��2����E쿻��h�΁m{۔��̹�!��Z��<�x����gEW'f��|�%��W.��m���\rg�z\����N�L���͘%e]��V���5��+Z�!�����HI�28`��� ��85-�ŗ7�����t��7/�z��9�Pay�j��� �~�%)����୺�)0�M�Y�m����r"j�ݿ�^���[��.�V��G:���U�'i��%��J
�)[$�b.� GqV蝴���Q�'P��.h���,��\z��y�Z#��?uɁe��qL���E��lB)�C���Ck3q���uOГx}�j�f�6ל����`��؆:�FJ �4�� 4;�o	*�t����?�-�ɍ>����c�-����	`���;�%��U#�t�� RM"��_�B��t5�.|_�fQ��֝d*�r�a�PT����YqNb�K��{�sUqȔQ�݂��P�Y�d�5�~���L�X��wnJt�>f�ĸk��L�v:Լ�i��I4W�-CF�@D/\��	ik]�U���E]�1*�-�[��!~ߦ�P�{fj�ZUe^��ȹb?cb�MH}�Q���.�;+���Q�� ��Oy��Y4p�U��\��Kp�����	/]�gf���\nuX_|lxf��LeA��~���	���|sQ	
��i�ɨ����|��S�]u�� �q�ݫ�@Q�#mM����u�������OE�b����V�1���30_X��Qw��lfɩv��wi;�<�nꀦ#�5���Np#;�X��L���<��{�M`���|���)�	ʡc6��h�j�40�6�SabXM�l���d��$vea�e-j�R�,HO�*Cz�%�L}j���X��+��U�i��i�4�{��P�N����l��C���I2=!g�����%��j��pTZs�ȭ���SW2 �	d�Y��;�h�"[�����*���������f�!��w�(ϸ��(U/��s�}*��{LT�*"������܀�찧�gWf�؛��OSi�5��d&�$�����٣������|�2�:t3-���'�y� Х���}T� ��w��ZLә��Lc�ۅ�;��<�Q_�tL�f��>�����]�$Ã�)d7�?W�I�mS��<�ha��pz�K��N!V�RR�dHΪ��_������4�P܈[�{M����~a.����T��Pj�]��k�>��VӬPWX� �3���]�8��6h����Q�a
[9%��ec.lz��`x���l������w�w���������Xf:�����\�}�nz�ǫ���F
��w�b[y�I���B�-�K;]R�b�7���7���^��D�����c�w%�=�:�C��
�_�'d?b&�4L_�'N��q�R�]Ւnϕ�FZS��Z� �G�������"f�F�(��EOs�K5�̆�e9�},	;�2�$F��0��,?�Y����UL��9��gk\�F�]߀{�����w)�'d!I���U�݋�>���9�Mm��?�סeg���V��ʂ�M�g�>6&	���T�_�Ѻרf���&l[�Ba-A7�)��_�E�.��U;�}�QG�}SK��%C������GJm��D���@�"�qH��Oi ��?I�����q�@ ��0%N����)�8�Ew���`�suK��h�p�P:.zo[1i~Ȼ���1�6�&G��x@�尩L=8�wR��tғ:�t6�E�=������k�ׯӈ=��11��	Y���r/ID^"�}A)B�o-�DьŨ�`�
���@}�䪦����C9T]��~�j��4Z� ���<�Y˥W��Ţ�u�
���HC&̶"��$�6��a�4��ktޯ��3��Dw�tF��9�Hk��� 
�cR;�ߘ�d�$j�x�0]������b��zTC�j��O^�
�N�$~]�)��M�rS���j�vC'�~N`���`k�WD�۳�s8q��4�R�'[�n�\<�-.(R%��#�x��5xb��-��Q���}%L���pF I���UH_7b�.�S	81i���
+��E��[U�����	��%�,�4Ipx�,���G�&��[��l.k T�-��j�I�[�Y����jQ���15\{����� �[^���㙢���#u�)���������4��V��L��*=ψ@�?�S����K�[����#N��@�cv�ޠo�1U���:i�G��]��g�>�;�rףڵ�4�'���0hU��{g�j�~����\���9p>!�!7��^`�P/��88���X�$"�� @b����緸�x��l��EJ8�����/J�vW~�7A��$����Ju�A!J�̖��g������k3��Z$��'��aǇ��hfR��֪J�/I�q�Cc�P�d�1��M�S��N}��0ʱ`���q�&XHr1��=g�K��������j��ڇF"`��nLo�EJ�A�sDW�'~���c����Ief�(+n�}�w!��b>�F>�'.��jݿ��z<`XS�<��m�su �5df��JQ��A϶4oG�4�2M�{7
�;�)d�GF�Q��<@�ڋ��Gsb'���~+��uk��t��
"�O|�}�� h�Mo��i�5����(�:�ۏz��|mR�cU�$n4,�'��S҄��C|A-��m��!��\���[J���<��?��"���j�ն-aƨU�#��[p�����RsЍ�đ��n����o��#���0����4P�۔5��?�&텷�I��b�v�Y#� �L���Ҽ��N�Te�nK�"�c�ΐ.�l�T�����G�-�DnxK#K)v�i�����������nG'�d¦ָ�:���9��]tD^���T��a%�l��aX�������G��w������϶�$ ���zD:�#@���p���E��LE!�����F  Y�މRq�22�\�u�0A��q�x���ؚ�" �I�.�5�t�D�{��s!�t�J��	Dec�BFF�����g`�Y���V?�4�{����E+��i_�T5������m��%��AE�C���l�9���s�3�w0])�GB0�Q0E�X���v�b��:���H� ���t�LO.^��&U�E[��O!n<@8�]�	9�(
g����fk� �U��\ώ�^k��"c&_S'�;�}Ģ�������P��5�X�D�Tct���pNgؔ��bJ��G:�����|u��6�A(T�[�1��(*��%j�{��iw�:�@zI����Q�csUDz+�h�\��UA��:�Zz<�D��Ժ�ws飝=��_�������gE&������{EL�9�����$����"����0�/�Gϔ;Xis�hN���_�d�Cr����~��[��"TQ&�7:�6uY��z�&x�7�pQƝ�8O�Qn�H��AkCϺ��4%i��Z����>������j�<g����,��.��ڡ���*	�ҨaaYa�&���S��0�'*�(��핋���j|�l��ZnV�=�������g�p7r�S�i8ߘ�x!C*�i0d��Z���"�ܣɲ��nuY�Y�Ü���y��Q~��ʓ��1��$J+*���L�|	�>z7�L�3A��r�a=�?L��:�F�m�`&ڈЉ?�,�s5��nP�E�^��w[ء�Ͽ<� �ti�R�e3��|��xyt�0y@BJ=���\M�p;��웻� _���󋅢P�6����J���ϻ<�a�;(���ٌg�b�<��gU�y����\$�+��fνP{c}�G�3�	D�����9wcN5U��rl��$��+��Ĩ�(��h\��_
ӹ�bS����p���ᳺ���ϨN�jG���2}MmBl���f����#��`�C�����IL�'�O@�|�cg��ȃ�'�@p�wD<n�k��َ�Ok ��3�������3�*���ХO��_��Br��/���Kd�/���#e1֖��n Q#��Rp�������)�xx,��+���B�L��&��0R���خ��5����I>~�����۶�?5y��5N��k��E1Pp^��@�k�8)��! �1�)�q���-;Q�ʝ�j'��r�4�;R���>�m����\o�k]q�]��I�.�kPqUf'>�<�&/j��lG�U��YZ�a� ���x� )�d�� �dY��䩘����t?��fl�7�� L�\�~�QQ��V�������"˔Ӿ郷�>�n�ja&5��!�SE���Y�KXj�9�I��iK|��C�A�U��A@�r� <�Q�1K&U
�fs �� N���Ǜe�1ԛ8���U7�έڿ�ɣ�n�r����@�}��$�`�A��A�e{O��b��D&g����(���^��2	�)����R=���(U�0��{s�:��nĂD�ِ%C������@>|����Й���bm�8)�[�uݮqP���Al���E�"�W�(Z������k
3/0�r�[D�B����ꦽ�u�>��~ZIꃘ�8MH�V�X���쎤��)4>�o�E�a�e�	r��R�b*R���"��ڦ Z�$����9����6�GE�������F�E���6u�2����?Km���]opb��xJ��ػ���MK���bT�mU�:S+�{�@I!"��f���;F�{�疊��C�����xJS��@xT�����n�!-�}啂or��W��=���V�d�G�1��^pug8��ZN�F�TP���-�U�V4���P{�I��o��,�or1�������d�����߇
�Β��Be��3�~P#��\T�ph��Y�����>Q�ԗ��4[�2�g�ΐ�3��;<}���n����GG�`�J���r��ff�M�# �1+�EwCԧ^�{D���	��E�y!)��x`�;/#�܍����:H�����$@*dy4.�Ԡ��7ԧ���e8~ +�`�Pn[|F~����j��}ᛁ���pH/��v1�uX�(��!vT��d�p��Ø�kQY��م����L��,������o���2�"��dn/񰉀�0.��p�(���t�R>���F��םs��N�?�tZ�7$�6���8Τ�UcHoٍ.�zGY;ak%����CI�)��"ey��u*\��K���`�Ҩ�Q)8$��3x��}&�@#����Z�u˷;<��;/�Hie�mG�	A=VQX39_^����7�Ǜ����:��df�mq���'9��(tn)oz�,�ʛ����f��	!�f��<W�Id���泔|i�����x�S��.��nsF��Nj�;n}�g�G?ͽ���2��d��؀Mk#x}�#����fF;߳���4�G㙎l�3ʒO�/ދo��E��SFwI"[�W�ObJ��Kr�,q� {� *G"�t�3���������d)���R�-���d��[���1�?�X����1�����A��F|T4����X��`��G,�Wn��C2�D�V��}Q�|�W�,M��)�'9�2�B�!ks/Q"�,�n)�oȭS�����`�y������h�y�|�qh���Ğ�acX������*VM��\F�m���S��_�IsiG��F�G���NXs�eҢ"���+��G8I�n7���t��N!Z(�w5��%�oP��Ug� ��r�>�b��=C����+�>�y��{p,��a �,y(J��i��0QF�<y���u��RG����c���f��g��N��`n��Q�>��H��H�3��>� �H�ʔds�:�GCܘ�J��1{�I��8�X���9��pU1yB��o��1Q q�Xk�-=4[�#�����OW`$8��q ��)� 0oሜ�˞�_�7���Z��ԍ����5x���g�@�ņ���K�O�a9�8(0��b� �%� ��~Qps���\^�(��c��r��
U!U^r&����(���ّ��>�� b�q���BF�2�R'��k� H���2�[BAgܧ�:2�ӡ��~�U�pEw���g�c�L��ܣ6E*ݕܿ�@��2K����m~w�*���+�����C[��'��Rox	*�0ci�� I������8�b�di��� m���Ty��R ��e�L����6����=z��;0��¯KB9)bU�Ÿ���
�=��S�S]�{U�I��1V7^����8<�3��j-�?�͜zߑu���n�Ђ�~S�V�w��o�;��������G�	�SP1��|�Ρ�h��s��I�n	��ڍ���Ny�<I�������#��V�j<�����V"�2�����;G�ę<}�T����B����ݒS�w�x� s��Z��al�Y��_{{A_bq����V�[�A�"�~�;&�N<��Z�ý��{���D�'�U"�X��y�r�s]b�/<�c�3�����S$�CL��Č��B�,S�=�͂����	
�!+
�I�|M�&8f�h�t��Oܝ~{��g^�"rL)��阄�KA�a�Q���R�Y�p�g��D�@����W��9�����{\�*����]։H�HΆ��)�,�u��6!D�ls�x�<?��Z|r��'�'ւ(�i���*E-N	.���-Hz�ߗ����cYV]�2���|ŷPZ�����$��3�|{g	_K' ���*/Vyt�4��5h��̀�Ӄ���� �"^j���4����K���!��aݱ�3Y]fO�S�8�1R�w&<�x"]n!�G���r�b�������Ud����_�(a�X���a����5��I[m����v[~u�2��mjx��Y}���f����z��7L}9s��6?a����{\M������w�c˾�L�B�j&�$���� ؉[�1�d5�Ǉ�+"���KP2`�~�N����Պg1]V���=�BY|�لK�µ�� E���
P�E�%��7U)���+�<���`b;ʓ	���f�����n$����xuϩ}��2��}9�\��UQ6����I�G㛩�\�����e��AP!O���}�/� �*a��ffZ=`J7�jt���Y�J�+����39JZ ����A��S��R��8@�C��_QH�i\����,�q)fq����#���-��Pxr<�A�/���E�O�G�\~,��2j��ezY��%2�8��]}�[C�/ϫ��!9����^=�5���F�i�;��u�e����xȻ73�N�p��Rj�/ה�t�N1}�J$�p
��,�j��"��_�-S�s�QSF�1?��[��xzo�iko}���{?�M��\"����Ǒ�7٬�{�_�sl���	�)�x��|�=I�ڡ��~�]g��ZJ{8���Qh��ۙɶ�g�`A|G5�h'�����_(W4Ff\�Q�+w�gÔi�K�
��5��X�tv�6��P���`Z�^g����?��T9�ϊ�o�[�1^���Ý�y5�����{�� L۷d�H�ֆT}B�֥s�>1����^�Bcّ���3�d�>���>pNb�Ѱ���Gܔ�m�s�PD�����i~,He��4d[a>�����(lO�:+���P�����~g)ָ������~.yR1��*V˒�$��!���u\@���ç��!.�ô�fM�ӈ�&��!�%�̗�O���(�;��%���By`�^6mh�oqzs%�B���mL;3~�o�l�S1"q��+l��*��ڥ��`��T�)w�+��/&W�Π3�/6�>9���&��W�#,>ݩdhJj/���Yd���!���t�>�8I�H�v�)��d��v2�d���]�[����oމ��lq��2q�S��|u�e����k���{<B���y靉}X龕�w�b����n|�2n�������O���y��B�kq�׼��(���8���ٺ���e��|�C�>�/9�)�L����3Fn�UJ0��'��yf� �Z:u$���>ř8fp5�^�{_70~���ń-�Fsu��byno�jO3���S��iA�++j�(o�,k%�K!�وI��T�����@Ğ]��o�P��5��I��^���h�hu�]e��� ���9=�w�����;>\�ew��TH�D��{��~�`����S�]�y���Jh�|�%Ԧ<���ߖ9{�
�L�qV��Ns�ly�gI{W��(*���'���G�L�bؗ�s�B}K����O̜���U|6�����0pGၿ>�ےF#K�*��͂n��Ӆ� L^��qf���'��u{k���M���h�љo�Џ�1�QTpp�lrƐ6�OϞ���fG~d��`ߤ��B�!i�4��c��P�b66D�1�|9���`�JB�C��X���z�e���uy>�V���3J:��Ԇ�����!X���H���rf,�^ʱ���[��9$��#��t]���"�c�6�h�:�rE72'JYi���8x�+&O���V�L53�݊�t��vG��E�7ˬ���FA�#G ��e�~53�<�)T�R��B�y����d�t������Eg�W~<zST�喅�D�i�Au�8�<����*g����9%ߌ�1QТ�f�\�4�]�D�9����4�3��\Y�^�)��\ˌ�������<�9_:���<�BK�P��7OL��'wo�B�����+�d�L�m���Ͽ'��d�'�f�,������5Z2r\}��y��g�����"�|!�g=���d�!��8L�^O3�%� ��fS��0ݏ��g�[�E<;ڮ�Kb�qI#b���@��'g^L*�G7s�A\����ڶ?C���=��vvEг�v����r>�w�R3!g
�^1��ײ/��r6
��T�ji�!�*��"Qk(m���c
�c-q��7L���I�_��~J��qi�y�������(ф���^�R8Q_M]�h�b+�=�TMO�D8��ί�»w�l<�Le�wP��;��U�O��1�w���Φ��4�刖Я'^��Ђ� �zp�Gq�9�~�����O��<��� ���v���u���Q���Cf���U�t����޷���<�`=�k�����K�E����x�sX�<b*���N��^f�$�
G<�E5�%�Va)��;����*������ͼ�)f�kCXCj=j�]<����5?��7�%���V���ft���Z��B���΁�u�1���]�B��Ӟ�W�/�}o5F�?G�ڢ���ٯ����c$~��j���yT����Ǥ�1�i��|�U���Q*yq�f�W���E�����D�L,�����YM�U{@�g���Ym��u��*���@�Q
P"�\b�4���|Z��r���%��9��[�Q�tS����srΧD��󀺌�ޡ��r�@���t3�9 <�����R����N�k�2\�=���`��R2ׄ+$*֝^�9�i�_���kn/���e���]�F]�P4&��78�t,�ZT�U��zv}�
ɶ5��{�ǹ�O�7s���=	?/��+�ݪ�O���W�@�����k�|��8#��H�5���񊲑�I�G��y�RT��X��K��[m��sS+��zaZ��.���xqR�^����\�9Ci�OJX�e�,c,Ts;���	Oz,U].�/�l,?�! �1SZT?dˡ��:?L�@�����c��b��.�0���=���a��68��E�I��n:J��=��@���Ln2�{��D�
�>^�����)�W��w���3ͩ_�`�<J���~X|w��M�#�<m��9�e�ҭ��$KJR��:� Z7Dڬ*��1[<�&Q�D�����Rʟ�"׸��f��_d�!P<^ *���`o�+��]Y��_͆��&�X�/ӥ����|�����	�ɩ��/-�en�dv��p�,�v�/_�Dw�W�'��E�g�I��E�Iwaz���}F%��������V���E��(YLfĤD�������Z�����@�Ɪ��-X�H�n��̰��&��$f�n%�EiN���JD��8���z��I��%$��������0��O�O񚅸;���bS)c���_w��ț8����Gw~t��o�l�ȍH�H��A�%�EWu�u�.|+�a�ׅ�ۆ?��䈈�l3ͩ�V[y	Goh��2t�*����ֿ�B����"*��N��D��N$��2��/j����E��f4d�w2�y�F�+�`�9��$�򤹌�ƕ);��@��i/3������T3.�Wa�Il�"�Kix� �zeV	//��\OCI��anF�v���(Y�J��$��`m�r4�ggr;~+��Ak_��l���t2�)E�I�V��'��zD|$���vEW�8��|V��u�TD
�����c)M�<��PN��n��1�<���!*pb�р���o��|�/������TIc���ڢ�Av�,�.�+>��r����)�q�ي�����W~v7�f��C�e�T���)< h[M4F�u��V}�jm)W��^0�Ab{G��>k_Q�wU�����^�b�N�6�C��:����"�2�a6�a!-����ϯ��:ii5U��Ÿ����n��IװrU�a9����Ft��ރ��u@3���t9��y�	��&�ɍd8���(��	��7!�躃o�@���]�}�aJ�"���̡�����{3>R9�4�F�/�p0p��l.�+���������@L�җ��w�/Đ��oO�)�C��Laz_W�R�/��rB)\�0D`�����X$7��� R��/[��8���P�ƛ��pF��p�"��:4J߽_.O$Tu[�O��r�CT��&�P����� �K�yl
kndЄ7���?}MhU��m�$U�DI��#�)@�;^%]�	䷹+MAx$���v���|�!3cyt�7KbHU��j��V�4Su7F��9X��6hX;�P���|��R�Ju�p�l"����lh�S��b��RD4�#,\�A3[��*��y��>ξ�d��f��{��Fh���)y��~3����w��>[t��Us'�&�s�a�^���uQ#�b�u6)͞�T4-�'R0�����[��da\�-xc�Z�Pg��D������	qX�.��j�FOH��eO�.��]��Q9���{Q�*�E��]�����df0Q�#���?��p�*v���!�����\�E��k���*�'^z�{�J�7��݁>��� � ȅr�7�ڎlzL�ϑd���_��A�c�د��YǛ\��`쭲U�^��2\�4y=�ڌ*O��2�Df�ޖ$,t�������,���yq1ͥ��]<�߉P�X�u�~CG�T�D��%��Xx��t��\DqꃳBǂ�ϓ���+Pr�����Q3}Ӄ�nkS'ԇ��灆�.� 8q��>�;��=?��Sq�����Ҩ�+`����rT7�8x�8��\,>"o�[�!�Mt7��#����W�o�x`a�"x�W�0�J��̏C�x�*���e4T�{-�n�y��y��QFGw�� >���E�8���a���z�syCw"�Z`��>��
�zG�c��}1y�m��54@�.Ǌ:���2/mp=u�/���Ff�ЮV�
���:�?���V����9����s��y�cNş���|�ȱE��G*fb�F������f�jzY���&y~7�{gx�(ᗤߧjM����$���3�d���HÑT�{�m�9��:齕ߗt����1I�K�CP�Y��+���;�W&IqW��x������:�L�����T�TF�)�р{�LXs�i�'��%Z	_�K�`��0��rBY%,��s�c���MX�4��y8��x��d06�[�����^�lXż�;���	 ˯�!�����Q��lR���Z3H4�ZDEsk��d6{�G�Itx"vtO��s¸�y����'e��. +�~�T��x�DTyG��%W�E�Y$��~j�CjI��b����S]q@����˿�qF����V��IԖ�lp�P����A]y\����]S�Qrm��j�1��Տ���]u�C0���Ŝ�dl;`Ba܊��&�]���L��� [����zU�����]5q����-.ϓ$���`J?�A�o7��@����ă���ŕ���et���r�PZ CH�s��F�K�-�����m��B���]�Uwt�lb�l�<�O7�L��·�`W[Œ���Q�n���	|����5����8u�]���r���OʊL���x��z/�%�8�ɷ����v$�21���<��t�xѾR�!��p�d���5��X<��%$���������������p9�Yt[��+M�e��5��duS�� ۹��/���D��j65t�;i��uA�ij����"B��gC^h�A�x��r�kj��D���KD#�l7A����?��	�o?N�*�r4q&��D����f$�QD�~��2��c]�Z��hp����nV�C�N:�7M�5�S���=!ma|��r=f�O��AP����8�y�P�t�8��)�i��(�6��.	�s���:��?��-?�e*[l����)S1�b�c1r�a	c��5�.u(��u�q-!,[��x���Q�Ķ��[�$�,-
��qO��FM�,=���a}��=�:�j���?_��U��;d��ES�)��2eHf�����'s�DT߽>���C�`j��L�d�l��'���"�����%Z]�LJI�)<$1*�����\���OK5a�@ƞ��W	''��O��c�#v���H�A�t�Av�%�l.#��c�/���j?�ȿ������δ��Q�돧��"��)�Oq��U�����s6���f�PVšK#����4��/������Iم���	aq����v��2
��XO}��VI�6�l�p�t��M�+U;�"�BݚΖ��A��-�C����L�r�i�˱|��zwNdU��X"U�	����Y>�K�CI���\��كjiQ_�sG�h�`�:��ǟWV(�����oeq��/qY�+�8��o5�j/��dk��nwZ�1Ql* PgU�����.�-�A����'9�yRH&�}�#�f��ؚ�*��ߓbZ� e���FO�c����{!�Fp1P�ģ#�����;7Zk���)�45#j�
og�?ʑ�J���{�R�u�%f������7���l$⥯�"Y#F���8���g(��)c5/��2���:��?k2�g�a� n�S�hG��f��|�����X�z�g)X˯i��/���RRg�z�%�Y���zO�$'��4�ͼ 	(I��^��L���3�Z��e�퇒�Ep}^�!��N�"��R���Hĥ�fi��ƫ�c"�2�oaāS�{s[J�$���(�#�ͫ�]�e��AW��}'0�x3W9�J����k/uy0��]��[��\p���~�P����	<�9�/$΋��?�IFL��B�|��h��9��jw��'�Ս��YŦ���X�粌ԣ��U08S�;$�C���4�jF���B>Aب�$��E�ò���a&EC����v���� 1�bo����f�~�I��)�o��H�i�K�΄��_�q�:�H��  ��T&�$6h-��ɽ���![��	��)���R�G��ꛈa	����E�Tۛ}���bH��`����	V-��A������~SN*���ݣa?0�(�V�$������.�~�5n�z��e�Z�x��e���B[�9Ϭ�m���"�&�K>��
F6Ͽ�!���RuXT���#x6���;��p5d���C.ŕ-S�Q�����)�g��W�����"������t��Y�� )s���2���,���y�l����$�Ud[`��oت�kU��d�~@<�=�h��Pz��R­^����d��qzQ�A�V:]L���5���u`.g�SPl�	_����@)���4:ց��+�R��5`����wmd$�ˮ��|@��L�ш�bl��&}��p}*��~��J$���:W�ꎂ
vH���@?R�~��$�j��Vd'D�;�����kvbR�<�Pc����-.R$��3����U�=)�{, �,���l䄛��VBB��l���	'�9}o�PsJ7��a�{�hـ�`ܶ��t#�����ϳҺ��SsڔH<>d<QP�����&ܔ�����Wk�Q�6�8����ў��NM�W�$�P���x�	�~�q\�X�����W����%`+i�H�I�0\���8꺆�~��C�!�z����nL?k�'��2��Vb�.����7�_����'�����н��A�%t��|{K yN��PD��|�xO6�	�Є���!��@3���,k�LWx�VEh\^�j��:e���5y�B�������6���$�������hbN�m���u��8D��M<�M.�T��� }~ȹ��l?����<x"b��ʼ���(C�9Ɵ�ql��=��~G�Gg�`��>]E��w{C�'�����2(�IVly���5��|,��TJ/�\A)/��J܂l3N���GOUdZS�V�4o��֖rX�Lk:���*'��M�r��-�<�O��*A+B4��/�],����t1�ٸ4��)tҳ�T	���ȇ�Vt�^�H^|��!o��2�vb���HL���hw�e!p����te��R^���~�N�dd ��ZO $��5�+V��a��mk\5W������9Wo�8�Nu� �p_���P��~���Pu��!6$����58��(4�Ȫ�D7M��V��\�'��h�jT���F� �К�>���U��	�_�4��f�b�������Ϥ�c�XAB �(���T�x��B�W �?�\p_}����>�����M,��oS�T��j)J���IJ/2� )�ӃH�~�����]�X�U=�ج��x���HZp�^�<tI����߲�%�X5� ����"��a�F{Yz���������]�!���e�Y&�I:`�_�f Hj��x>�����x�jy��!&`��BɠXQ�
f�`]��A�_d;x�:Ik��K)Ǻ�A�gA���,!q�nI�ņ���;��B%��k�OD�h-zA�f�(�:)�I�<� Eϼ�O�!��S�6&x}c�ܯ��Z�� $u+8����]@&�`Л�z��[���B�]Jaf���[��n�h�M�%<��U�c\}��t���V�ϴn�s%���O���ˍ#mQ�iɩV]+~|�W�����%}���&��h��[����Q:aS��]���
J,�.��O��A�/v���/4��*m/�8;�M3v������@�i����A+{�?-�w�Oo�άR���bT�!�`�HU�-��LtBy�D[��r�{u�d&�d�c�h��x�]b��A+l�q�RBDÖ2<�_~{��J(1{�W.�5}��I�6� ����~,rX��w��ݪ?}}a��ۮ�6� ���-��&�l~}��������D��--�����z�Q� ��^_(��W��G��G�{�����V�@1�H������A�y�֊i�G��Rr?zt����6a�Y�oa���c3Vp��z�����N��
na�J���nk��V�}�''P�[��͏':t�� ��z���켓e�=�Q�Rh&>�Dp�W<����Ѭ�C�C��ɍ���=!M*���>g�N��m�so�.^'C|񞊘�m�n�-_w�bT�lni���[�ǈge8k�󣸸��ȩ� jҁ��;=�ђ	��[L��W?�[��p�%߄Ϭ'%�.�"�L��gkk�>���xWØO+}��X�؈y��a�������~Q����.����c�\��7��}�F�=my���MK'h/Y��}X�Hjm�M���e78���V�G�<�V��)	�Q�Z���!(��7G���C�kH�+�u�lI�Rr�V6S_���+�j�G�ˑu�w�� X�n���%�E�>Nz�×�:LJ��l�F~Q'�*ɇYv=D3�8� +I�Q�P���*k*�_��㹴^aFT�8����1�u=�9E�����E�
�=���S�P`���2R���� �;� ���<P�K�Ѝ�~�	�0��4�J�K=����[��~�bBH����z��O=������\���RZ}��W
P�j�����}���2ɸ�����Þu�6�]��p��5M��̻�ht��b$紼B&EU��t��b� ��<���;fO��Ȅ�Bpd�~%ƨ��wP�7�d�E�;;��%'�v/��A�*�Ό�CD��7�K0���V`EǑ��'����:k�6�G�2'˸��ZH���]�Oa��J�S=���ު�ߗ��PNP���"_��%9LRt?���]�~?��6�!�m� 1:�)�sM;��ȕ��_C�#�XF����h9�^��gqFiꡒ�bq�u��K����4�� �w��	V�`'UX���^�_��q��hb';�Nĳ-`������%>y��"'�a�K��G�x�bc5�I�q�`C�����1��-�O�ݱG	�����DQ)��!4��AH�������f����>�v�]�C>}��:g����Ka��K��n��������NnMb:-�F��nT:�s��t ��wҗűM��ie���7�$ڗ��OF��2c(��h?Ӛ(���j��k���_�h����[��n���Z_�^h)އ����������߼���`_��eOŏ�1_i�'	�]S*��vJʷ��n�������̘�Mļ,��Z���[�mu��V���Lk���O�V���e^sWp��[(T��q� ܃+���`G��S\݃�w��k:�X:��~L�w*$Ib`�/ϩ�����8��%� nԇȶT�X�'W���u��$�ˢ/%絍��KK��/�)�Ҳ�Aȩ���
7tw�8�rs�B�4��0�u���1��`�l?|-2h;!�]E�`�0�^Dj��,.w��C��a����,uT ���A��}���eQL�J�F�4�����H���8��> ��.��|M�yl�,J���
�os������#�>
*�}j\4-_����"��UhMj��t�x�����ޯ_W\wT���yTaxX���@������Є�9yH�7�W�h�M�
%mv wa�X���@&�����<��~��3��4�W�]*M�䊈�F�����~<Ő���W�⃫HT(k/��W�pl��7y��_���Q����B"
�����(؋tϪ3b�_x����]��Έb/����Ww�s-i~;�!�JF���=F	��J*!wb:�\����t.�=�e�Y�A�_r{~$���*�����ܜ]-��wZ_��o��25r�GZ�hb3�Lr. 5z�9��*Z��&�4���tL��އ5B�����Q.�@Y�&}�\��РU�:�����k��}�����fl%���R%Mh��4�dAR~Te�N��?b�����G���k_rw)HD
<�p��wh���´,�p󂗒�h��#����Gd#PZw"]�Fzw[J�U�`�'s"s76p&�C,��i���s.ݡ<���{���"�o��0H+�P�*4R����BM
���J�$A�'��h����/�hd����7���>��ZLhY�Ć,�X�Z�h!G��Ǣ��v
�|p�FS�
|�&/���7w>3`a���@��U���P�ng��<f���DEiչ\c׮.��}�n����M�ţ�܍�B�?/����Y�@p������s��-}��F�)� �����h`�U��@��`�ʬ���ǵ��ԏ*t�5�d�=��/-����O����l�F�=�A�g�G	\�n��<J�~�Ãg�oi�y�� %�75�M�f"�3/�6��}���i��4�	t��� �vs�K�����߲?,��<�1��BY��n4R���e�?�kx������C�v�)?� Vf��!#��~nA���]ܷJ[c�Ĭ�B�8GDF��~K0�Guw�`\������KD�5�a���,Z��+�X֑Z�꠯	>������_��m��E>_�϶7�[�h2�C�&	q
�6����G�r� :��.���(���xs�׏m�C�v��x+�,��k4ۄ⥶�gh�D�Ǭ�q�p��$iS��I���&�%�@���7r ���CAh?}�T����kŰ�(�]l�J�����\/�+��� ��3z�Ҋ���~Q��AS�)�S�ОŹ�?\Ƞ�NJ���Yt���"�Þp��㏀,@a����rO����z�C�la�7|̈́6l��X���S���y���WEO�ݮ�-A��@������9���%�О��n�����?3�x��I^ �)��ٵ�=���845�a�45E+"ϝqD��s=;�e�*I+����\	�S{+K�˨�v��֗�~���!N�"��^M���00ųG�}���88��7yw����+,XI�˲EB(�F�P��ΐ��z�P7A\�y��g�t�V��͐��4ɂͯ��<�X<�� ��u�~1l%H��9�N�рW�����_�>7�ё�F�^ݒ����~*(��s���G*z�������;+��d����H�u��xDZ�<����]Zs�lП��a쳽����@�e{н�X]<;�؏��X�)�� ���|@mY��uv-����b?���A�-��;����N1���#Tt��5-K8C���n8�G������c��� ��x�7=�������%�|�g\��\>��	B�3��;]"%�~�!w�mgwPz����b�+=C�A�t�X 
y��4`O<�#[� ���ef���$ͯϓ�p\sxS.ds�v[{���d����廘 ������%m�E,�v��s�����+h����{vAbSEI f��$[��_9�:���i�@�ϡ�[w�a�纠^���w
fc���?�B�@Y(��9�`vQП6M�9�>M����:���4����W-~�D� >魶��y%,!�HM[O�6���$q���#^�]��G�ɭ&�����.�m��!�m6k��6Q�` �Ԫ�ZL�X�e,��'۲H��0E�h$\zx��̞��@n�
l�"9�+FX��� K������/�h߱�B��:*E�4B�ه��ߖ �����!��j4Q�j���ЖBk�;�H���t@��Q�Pr:�|����#����\S�qK�K��q�����y�D�Y ~��F*.ٙۂ�x6Y��Q��J��5��28�(��� �p����7E�if���RM����x���3重��tSd?_(��T>��f�C	du�R%[w�ڒ���1R؍�(ϻ�)�<q7Hk��Er��ǆ�	����]V�2�}�[3ΰ�?��m�B2O�¿m}����yU������u�@�e|�5S\�|��D�l�V��cM���KT�����#�<ϰrl�Uk{77���O�9��2�i����9���U�K�]y�b_�[P��9�[|S> �8����O7���< �=��ZX��VT<<qB���j̲S�O7H���_�\��i>�|��k��8Y�H�:���Y�K+c5�ڎ"�_@�9�}5� u�])���/.��Ք��A���v"����}�gVˊY�	�3�N{��r�"�Џ�/��WJp�fJ1�'� �"[UXb��fVNKRr)]	��uqVZ	H	/?Vz��yt�ύk"�$��|�+�6p4��+�Կ�#�£}���E���б�-����T�����C��/�z3~�}�h^�5m�� k Z���Țx��{&M�lԗ���3Aa��Ã�K��'�ZK��2TȚ<��>5{��h����<��ec��.��ԢFw��ca�Z�K����C�`�B�%��\�M��Z'����RҦ����eQ� �}g�����B�=jh����d�G�?YQ�5�j�/�5�d���>y�Ļ~��� �6:8u���Z	�+��
ߐ���\�r�X��Xx��������Gg������T�2SC}�Pfa�������@�~0����Y2X���ܡr��X6�=W^�����[�;���w�z/���SIa�Rvꪾ��u�H�z;s���V ��˶=ө��&��U��fP-l:B�zk��H��u��X<����u�N�@���Tȹ��8(axd�=��]�f"S����j+��o��9z�����u8�y�V#��w/�Ի�� JxbG���|� @��o���\�ɷ�h�f!���zT�`O�^�]�1�&�˱�@n��q'X����D�Nѓ&�$�=5��'�O�A�V�DAg��@*F?�Q�#
^����!�2�(��(@)��G�*.Bc �̺��c��u���8���/��|@l�Ot��!���I�Q��E���)�V�[�f�+��:5�XP۾K0���v>4�|�1}p&�pԅ��\�O���?><�&�eQ�=�=��,3��	�A)F!����r��
x@�\��(�=��|7�UָT&[��T{�§vuD�� &O*�t��$�2s�UH��X[�%�	��.f��re�P>U��g��1> �q