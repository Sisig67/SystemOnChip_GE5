��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����� ����m��Q�D{S���;��ie�9ߧ)������o�A�o:qlQ�����!-�k �|�ʯ�I�gr��A�PmY3t�}��`%^�"��/A@5Yϧ�a?�8��*���p�1/�XSL(����;1fKv���:�N�烋�������}
����~"�ExW�mS�p�$n���MB�X���dLqp�r¤1]��1NO��	���Ǟ�{�����A>���CFĈ���l�TI"I�Hb��Kh�]�����	��Q�����Z�[�j���֯���Mv�Lr Ot��(�R_���,š*Ld(@�v�4���#A��3��S��V3���[��Y"~{�d;(��='R�Ğ�.u�LDV����]��fok�x���琀�C,L9n
�}�q�d&�h�͝T��Ee�^�k��F6 �c?��e���FL��MȤ��iu���
3栍���m��]bM|�(.��yD@�PJv�g�D����ms'F� ,�MӰ��X��Y1� ����X֛�,A�&a=�*��u;��S������$���x�E��0�����v��70��m��H^��\kV��V�v7���i�,M�V#��w߼����g� TLY(��f�@���(���Q��D��m��;��l����B�5�z�L����w��#�����?�z�/$̲`*^�	�si@�q�3�9��y���=I��!A�*iR��Pr�R�.���:�L�͠�$SF��Q��ۯ!��F���u�f���k��݀1�P�(��b��ݘ�y����<�4}��yJ7��s;�n��t�[�y� �\�pW�݁8��_��8��w����q��#ZC��6��ީ�*SJ���PC{W�7(7�>�����[ 1�ۺ)���t�.��ǝ{uj�J�-+���T�x�f����G^0P'��F}��gD
w�:~�AvY�<���?�쥳yЀwQ�~.�Eۖu����A�I."f�F4�������1��R3=eۙ1�"�p�S��:K_"�9>P3��i<���	q1Ka
���4]b�����v�3Pmm>�Z׫����}��-Y��^y�j�0B���m�Yx���������I٠f )v�� W�q7�Y��xǸp4EW�7:��RF~��D7�V�L�&���cjB��0甅��;=�g�ْ�:?��ER�E6a���F����ZMa`	9'�]h���I*��h8��t+�g0��l�D�\vo�"8!ll�WM��v8`hi�?O(+uOA��%���mCy}���,l%��d
S��p�p{Md�"���*���ԖÑ�m�����4
p3��ک�Q�����v��КS^�F�.��7g��J���|�����ބ���'���g������{v��ǧ�<-}s���rK�؝�q��u>P��?)��`5�Q�-J�8q�v�y�?m�Of+:��?�7 &E=��О�s�N>A��2���ܕ�\ -o��l��m\��QG�'��s�
q��J"F��݂�B9���6)*x����� {gRs�cҥU<!�����;����������%���:x�,�8�o���qu���^䚥��0�a"���3���Bd�bN_����FU�(��d�~1 Ǔ: ��ᏐR�p�H����U���`������j�B/�7^ѫ���J Ukw��G�`��B%;�<���$(���[�X:t�k�@r����ZU9�ݭ@e�����(�'5�E�p+g��I�������������;Zi_��2[^ITi���� Qm����`b�vE��������s�?��b��ߏ���xظ�m�?����<��*�U�\���*�PV��l�y+jS!4o��Y����\a���ݥ�]BIθ�*��k4�S���;<�lY����³
q����좨���䓳�
���=��ՙV�^0AcP]a���  �с��R>��u��|�Z�,�:��q�#ݶ^Z��qM��!������!;sE��?HWVxUK-���r�t�x7vy������WP�W���[��r( �K:��r'���-Քp��Y�t<k�g|Օ��aʀ����H�%��V�R�v�eD;W�c����a�d~�'�C�S!#�)c���ԋ_�VŒ:�	N_[D��@�ͥC�	HD��n��4"��o��"ګu��ޅ0�$ɝ�U��\�s���O�0��+����&{�W5P�3��q�=�+&��|ZHb�E�$�-�V]���-u�!��}�*���4�R��w�`�/Uv�Rw���D���e�����3�*� E�Õ�黏d�nS�o�h�nǂ�Z�]d��4��26
s�,��is���������O��):u�x5�9�np�Wb�ߍk�`�t\҉�ɺ>�k�;�W	��-u[�|�W~	�����z��ڱ���_�s�I76w�g�Z(n�fw��u��b<M����[��'��vH9�j��
���`Z��,��*[���:�f��c�Qs�+ ������"� g.�w��-�H��:jt�GV/��3��S�
���R9U���8�;�b���ʄ`({�O̱�5N�S��ؓ[�X��v�4����Oׅ�ؽU/�3�e��_��F��B7A�Zއ�!�޸,e8;KڔA@����DP��1����ª�P��
;��G�	�Y�L�Q��d(��,K�&������t����X�˕ӱe����E~�wU��hk+�`�7�l=�,u
m�@�z��Xؖ�j�ӔW>�u �qD�j������x�d,ö�w}dX�h	Hy�ֲ���O�(����;.��~e<�t�FN�%�AF�/dS�k�t�VBG,��+X�hPZڭgFzHZ��[�`[Y$�����'!4�	g��}�>��ؠ]��%"AYq^�iO# K�[�4�N���_���GzM/>���!hI�s��S����|�?l��).����|�����0GI=Q�+rd#�C�}i@"ݓH=M�he�΅���S��CxAJ���X�".c³]r�������D��XE���o������}�	�⁞^W�e��$1z�7�GYM �A��������9��G��CH���Z�LD֬Q6rK/ׄ��{%H�v]��<��ѝ�ģ.RNVI��w��N��ǵ�ye�6F��^��o�
���V�ZP���_b#�y��v=�]�V߀K������\K���-�6�Q*��Iw��j�W%P-��6H�f�j(�6�$���.��d�?'�������6��t"s��CQ���
t��-�Ӽ	�t%��N跉����Z�ɫ�@�忯a���J�����r�3S��Z�:�L�/�H�;DB=o����]1X�FՑ��Ip��N'�
�N
�U�p�M|[��}�_�F��^�Ǆx�����W���O�I �n���n���.JQ��"���c�:�Dvu-œ-�$-�ĩ��J �C�W�SF��k=��ʟ�������������  6����=�p����՜_Ah��Y:s�r�
����*����V��
����(&W��SO4(g�cQ�e �S!u�?��4�Kp�7��_c���� �|tc�����xH'�m}P�MS^��[������(�n@�wH�=,S����hWO#%b�\����I��[�:�����=|�qv�xT���&�E��=Um�H�6/����S�K$�$���v]�
m�t�F�:�?�AJ���ET锽%8n��bpS��D��|Ǹ|k'�nIm�p�j��P���*��"�@௩V��R�i���`��S��;�Η�}#˕w-�F����Sk�ʝ������DGXj0&����f5�c�q�w�	�$+�]1@���|)� [T9�2�V�1q6�+'a��m�,�Z����'9q6=ǒ�<�N4԰���l���gCC�-���&��6I3_C!�gf ������#��5���b#}��.��N=[�����1K~�1��R������=�����@N9!%�#0�_2o�s��o�7�ae�U'Ho_��p�9����i�O"���tdyTQ
v�����<���n��ا�zc_�Oa]�zk Ww��}6����g�PX�4�B(���V.�Y^ʹ��ÿIZ�0�qT���PM^�(�j�����0z���j��S�ю"�7�h!����d���p\�8.La�ֆ�4_\i�P@�ߋ����e�X���֘�{�y�t��P�u l N����|��Jɻэ�+*Z��>+�]�]\ZV��ϡv8���)v�j�Sކ�'FY����s��h$�f?j�uH�F{�4�>��3�������N�q7Ѵ��3�'֟�*�O�}3=(�{��L�o�Q�e���|�ڨ\(�C��?��+5�Xҟ ��~���nCTYLͳ��{��>���*�jC�5�}g՛^C
qj�6���sx��"Y3#_�K�te���o�̀�t����x�����Ӕ�"z��u��*�w�}�&E$���9Qb��c������칪;q�z:��6Ղ��&�CSW/�ڰ��,9� %�uj}�3Z>g��u�י4l�zf�k�V���T�y�����r�+#���UW��l�&v��.>�&˷�ߩ���q�L���[�`>�ɵ�7��觬SK�O)�
��!��m
�u�eP��y-s����ލkGCRR��`�vD�L�Џ���Sqj5�P7�:��7'I�1�i�L_߉�uL��5e�*~�g!�;��zF�z��,F���-�i�c���g���DVQ��_5�#[���H��(��P.#z9���4Y��b�Y K�ҢJ=�_ ��/�7������{��[�5�׹��3oO�S�_���Թ��9Ej�7���]�#^��f�R N�ꎔ�7{�^�Y#�	8�z`CgR����G|��pOY�06�>J�:���N�&�,~p��k��g��ռ�Y'��H�U�~�� �G�6[r�U��B�L�W�d'��Fa$�%����w�e�0bsp2j1���b��2B���֭��!��	���bj����N�sD��Vy�D�{��~��t�1[u��B���)���_:��d���.[zx�9�& 7KC�Aǰ�𿶌-ՆAHB��ҡK��aR��݀`on�A-���f��������@^�(g�E�s�)S���ΆN�X��}��Q�[� ��Ί��ӗQYM59�f��������joY�_�~�c�b�� �;݁�ռ��v���],���}�"�+
���ۯ��/�n\&�T|��!�]L����\���}Jp��~:G#"j�����F�[�-(���Q�RI(e/ұ{�2��0�XEk��4�`��k��(�0���~h �$�/��CxI[@�Mֶ4U�WE���s�}��Ys�
c!t�ܾ�#'��� �*�	�ǷD>B<02ͽQ��
����n+V�ʖ���dqI����G�n������)G��w-e�*���$�h2|^��!gZ��W̃��Yt�z��CO&L�+�u����v�0�f�sI��%���ļ������H�8cZĭ�ɟ�ķ��h]��a\�Ҁ`%��Z���x�Ӿ�@��֧��ײى���r��p�f4c]H�tW�w�Z6ߴݯ��v�?yW��.%�7B-L�陮�7fAb�*����yWۜ��РKw.���_��43t�'}E�X��bmNWM���=�� RK4�h�-�/��&֓���u?S�+�b��~ZoA��<���F<�b(��6r�xml�1]�����K
U|8��!L66�XB-.�1Tc^�ݗE��nf>�5�����$�0���w(��#��N} ��"�?�bI{�>7"�,��0�g��Dۭ��D��H�}���z���b�/vh>��GQ�D�:АM�=>�o��9a��*�  �@����գ����SM�"�њ�Fİ�d���WD��G|�L5А�F�z9b��;�ﳩ��c��s�DJ�������V�9���ߑa��!Q����\[��Q���ߨʙ(�>h}+�A9�Ӽ25I=��)��,*N6�]��P�L���h[�𰺷
��N�`+���Lx��);�f���ϣ��߱�RO?�G�թ��_X�o�a^��}����̸__F\~?�B�B͠� ��Ksa�Dz@F����l���\3/-:*��|o�� �h�5�ub��.���%OY;Ty�/�U/`n%Î z��neɇ�B���g����iHʮ�y0Pe�L���]���rnS���v}%���9�h�{7��@�zD_�,M�^(���.�	���o@2%c9��t4���Ƴd�.L�{ݮey��V��,"��~�Y�YZB�b �l��Q�*��9�����t�-�4 �ۗ�q�y��?���?�
&B9tl۔���S7B�^�V;%7�
��옆I2����3�䄳_�ه;�R騮|�fX�n�0�n%,/�H�sC��H�`�s�D��Os��'�ϳ:�.���	�Ō[��C�5�h�E�{;$U��܌�F^�S���vq�ۂ����&uf��b��*��`e�K�t��}^��,��j$[����@_D}�(Æ&�W����.@h� .3��/���3Y����節�p�D	�D��7r�:�c�+��p���b��^΀��Y���*�j�Z�xO����+b��|-���5UjŃ��}?�2���ɮ;���Z����.��H�3b�B2\d޵�J.�_0A�2����wt�R��)���i��u�Ñ��3g1*'J�.,m�D���E2<O�Ni/q��/��!�� ���^ʑ�@�9z�N��7�w8�;�e"���I�cA7h$Y\�#Rv~!�|W�V���vpr���{V!A�E8!'�^~!�
a��,��9�����څm��=lL��Z^��2�^�_1��mQ@���������V��M�O/��.��2�����9��P�{%�f|�D(��,a^z�4&54�j�2�uU��t��.Ǧ6��3�ݲ���R9���d|}OxތꁚԨ�F�n�[��jS�;�k�9�R�|jY�d��_3Ж�蝓UJ��#��_���п�NEX�AUw������>
���L�*+l�(b٫�x��/���� �HAW��J�R6΄�ǩL�e��~�T7���y6i���{_�I��e�(X�3*IߝU:�0�;>�3E
�쒥+Z�{��?$r��kQ?�[0q9_�ߕb�8bR].�s���Rk"1%�����E�Q��]8e�wQ��K��0�z,K2�*L���禆c�s�H��¦
.?���D�������J��8��)�j�EM�=����<���Ӏ����=��hou���?��*��hP��태��ȝ[��["��*�����J��tUK�t�2(��M�"�Yn��yk+�䉏Å:e�M���{n��x�B���4~Ӳ�V٠tȥY>�lC"���&}�t��0���3��̃R�(d8��!<��_��D�J�Э6-'�����QsZ�2�����7�_�yAp�5��RI����>d�pI!���$Y��-��AY���6V鍔kB�A�^�<Dw��˭� ���AY�"���]��&Y�k�V�ma�t�RlոX�뵎;(װ�H��%��LgL~F�v���Փ�� �xg���s��:���	f�k�啤�D'8с�~�u� ��@��1�kh�Ftڟ� ܘA䳞s�� �t]-�`�'�Kj�[c��B�h`���.���_T%��
	.f�:�����?7Bb"�������?��/��ə[`4��B7:�Le��h����ŰZ ;_z(�Co��귶_V�^��^T���hu"��p�D��ō�9z0�� gI���x�d����hX�س3����������ĳ�����\�p�s��_��A��zF�@�1��To�A&	'NŁ
�u֥1��N�5m�����A9';�H>���g���j���L�,�X�1[���:d�m��w$%(���$ϧϵ+����z��ۯ5ƪ��\\��.��HY
�cp�sT�o�/�6L���-�܎K��[��ͦ����,gU���Uۇ�z�z�q�k-ei��p����� f��ݻ�Z���Z���!R�Qێ�2-zd�{
��3�u�����'����4�1��,�0�� Z��F�%6�J�2E��69[�#Exw��R,��@��B Fb��b�p�_-��	�$�Ȣ�m�.�%z�yvSJi����3m��।{1��Pά;�a��'F_YNT&Fߐ�ZdEo�����nu���v�eÖqmR�$=��V�T�����iKХx�3���vJ��g仸�9'�c)�K�6��Q������k;�@�ohz�q�토���"��M2�s�;����Ilz��L֨s��!>��L�\4�cِ0%SY_Ӧ*sr~�L>���T~~�V~epZn������A�(����ai=ˏ/'�c���0�T�ٟ�:}Ha���U		VtM%�(/u-N�iZ˸�A�C���l���[�����(,���>��+���6ƨ�dvK�T�<�x����S��3k�W,��{4t�y.��bͲ���G��o�ǩ��e5#��1F�	���� T �#u�s?��~���@�'��m�r�x�j%X���ETr=� }�w�Tw���22
r�F@`�gJw+c8�ޱ)H <R`�PHA4��h*���Z6=��w�<F�Ce�Əp\x/3�]�$͖���r��r����`=֋"��Y���0_�$;y�ٿ��.���:v�m���a�PB�Xe�?����S!���H�F=B���:e4�dWTF��7ݫ��H��UGޔ����9N��H��"�����ɴ��,���&���-N�6�E�d�!\�s�'<���n�Tǟ��)r��}�!�I��|?p�*��!���r�)���p�J,�)���f���҄����Tl4�p�in�"z��!ћv���<^�P��������xp�{ Ouc��7��ck��x�^�l�]߈�֧a,#��$S��!�ŋkX� l$?���p���L7�������$�@߈�/7Z��0������h�W1e��4=\~H���ﴧ@Ю,�\�ԅ*�9�|�h�Q�[�"8��dM��a�JEޝ'S��e��P��/`�u5��%<�ȶP�S�	�ٝ|��qS��(Z��\P�Wl�2������N@�-ͅKp�.���C�������f��r����3��]�0T�s������)�]�0	��8�I��5�1oJw ,��m<�
4]�
��
S�q (�AF�W��PX�o�=%ð�i��Ý��(h�Rq�f�FZkw~?z��:����$��.ER�����j�
�sp���M�5���G����Jf�����y�XGm����H���|l��
�����\��΂���5Crd|�c��%�hQ�~�z9p��N��!�'�bnQ*�;,�Q<������c���-�w1E;?��B#�L���'q�T$&�a�̮01��;�.ߨ��ޜ�͡C��1�=J�f���h=��s4	�NK���|��U�f/ҸVܧxM�
��ɢ����RP�7¬��x@�2�����_i����Y�̸�\q
���j�\�e݃J�"�9��)�(k�sQ[���NS��S����ٶ@�D��#/�
7}��?�W]���uk�\gm=9�o��1-������Ú��h��1�k��ed�w�N-}�p��m�iG݌�@B���{@;[P�+�m�L
��AR����Q�-k��R�'�nYH��
Ɉ��,�/��hV�-�����e����� �'>?.)-���8��?�u��[�,�Q\����,6�|i�8��*�}��)-[IY,봛�˳�̏=³iu4`��*����L���@r&Q�g�����2����Z�W�0/<4u����R3��N�)��.��"j�R��&�8+օUP�B����*v!_�a���.�� B5��־ғ#���|�	tYp3ә�4�@~������td��*�e�30����z�#�D{����ZR+垉���դ� �Gw�<�� �x�n�K� ���9�^낣��\�M� u�"��J�>��gt4�qx�ǿ��<����Ƽ�:+jsW�o%8��a��C�#�*���׵�Г���S��.Ed.�T;�D�C$?�����h{��\P��� �����K�B ߦ0(�bugĬ�L�ܜ�j��;1օ����	�'��ո�*�̧�<��J�90'������<ɱ����L���-�V,�p�v��I�r��I���������H�&J��=4��7U���3�$h0�r�g��עpx;�0�S�6�R!o�>W9���/f�o��i��&����O�hR��	�a��#Z}3ٜ�L:r�|�/['h�}��7/gy����Dڹ���q+��tX�Tt�.=��#M���%��)��l�
��7�B,�uT��>�ŷ�n((��Kbc��K-԰"Ȏ�ws�X^W���8�>���A�0�2J��
k�8p�"�ӯ�W��b�вN@	a>�� �G��iv��`���n[��α���1A���C&�oϛ~����U������A��/0.���L;��Q�[f��s[�<50�Ä�����0�� �I��.�H�OGo�z��|a��^p#3 w~Ѣ�󱡓Ba�Wz�WIs+��M @r��n!qEdm���(
�0�����l��xk'/�#,�� \k­�X ���d��V�4��{���q�Z�̹���nʊ��B[��>�����@�o�}��b�˱Gt�i�g�G=�(�˭��u� c���{��xa������]�{�zSNo��H��u3+�o���1��'�����_s��9yVĊK���FsZ�Lp���s�b�)g�&Q��@�>6�c =͊Yq��M��%�?x���_��d�Kb��䳈�ϊ���=�l��fb����P�S XC���C����ΰ�ط��nb�{��`R����w:�#k7���� ����+�� �����ڔ�� \F�IɆ�\��J0|>�L+������+��G�-ʨ��5�i]l_9|�*����/Ǹ��� 0����x�x���a�O���0�֐X6������6o����-�a�\�O�����$y�7G�	�An'#pɩO�H�4r��Bm�V�l�Ay+p��M�ߗᷩ����i��7>�wM�6X�I���C�x�ŽJ`Ԍ ݥK�o�܋r%?���?�,�����ɫ���Wrz?+�3#���n��#�Y�]�k�Ų����%��wZ�r��B��`^���t�O8:gfV2l`���I3iK���M6@���>uRL��0�i5<����?(ѻpQ�/t9O�Q^E��0��p+��X�H�X[�͋�V��4n
ؘ#�21�\�����_!D�1u�^M�����i�����WuW�%�&ϯ<��+&8��,��3��A�dw�.�fv�{��D�p�w:�ÿ�'T�{"H~�X��Hl�).��n�~L\h�i�ȸ��
D��`$���t�3�S�����q?I{p��v8�@g�}�^��.7�z�6{~��'�&U�25�+V���i��Vec�eX%�l9,՗`��Ӊ�I��x��P��W�V1�5r+֤+�І�܈��(/�+��O1�\�e�� �ܤ��%��?>�yp��;H40c�F#����h֧p>�\�����OR#C7F���A��E썌��Sj���=JB�qFJ��. ��b[{	J6(��C��~W���O�1{
/��X���m���ӊ@�p�%N[���N^�mLW |a����=쬨^ߜ��HZ���&���
���W�%����q��JR�����S���I&�I" �
��;i���۰Z���'N�x��5$���|�G�vg���8� �t9��|c�z��	�>b(��r�~3����h^G����-�ѹ�"��T�_��K����Q*� eOIg�7���B/8��|���#Ƿ>u̿��Yi�hU[��mc^�,n�z�w��~�\��������/��t���9� �P.&i*Đ9�җ�+9OLb����2#5XHF�ܧ����,>�h5��ܐ	OW`���kns�s?��������c��l ��AI���<�^����$e��Vd�~z��Fx�1x?�2���ìXI��"I)vY�\�^	AF�ݽ��3Hk���Q�x��wV�t�V�Jk&tbE�	{�C��7�b�:\g؇��QL&	�V���U�V�W�k�~���z���y�a��ؼ*��J>�+���M���nݵ�\��/����z�@U��{`�+ڵ��7@D#ԞH�Z����ﰛC�h/�⽥c��7�˽s?ܨ]�y��U �F�a�e�G�x��&k����Dv�k��K��~���W�Y|�Up�u�Iޛvބ�GiADk��XnNڃ5M+��r ��l�5�&.��d.&�Z�!�k����ў���J�Y@!��V8���c_�}����B��`h��wv��_�@}`�����z��i=��FD)r�0���k��:�����BDx;ojM�����u�z��tٛV����C/.�)@w�N���={Ѝ&�h�dݹ���U^vۺ��B�S>�
D�?�2b���b�y��NK|��m	;��H&k��.��nq��W����V���u#ҿ]�F�O=!:�G��KS�3���-�,Go�4���ˤ�Hh����3gm��U�@�z5���x����~��x#�9[�����VM��'m�v����B
�����?EM��En�ݒ���@0�f����Bi�$�J�l-+��>��%�շ"P���@l6S�
�� (D�7�_z/B���}v!��99}�뉂@���s�T�M36_1'I6���9k��`lٻ����9�5ocC��.�>E��Bm��H��}��E�F?\�PT<DT�խI�{��'��Q�p��څS����:��]�[�N�3�En2���Z����Z��6h�;Z�Z�:��P�V�����@�J��:����p�:ʂ��ȰMJ���h�5���j�@:�aA����b쒢{��myu��-����ET�m6�\dl�X�kye�ò�-�*�VR>�����2cx��� 
�MxЈJ�FHX['_�>�K�L �)��ڎun��9{��fՆ�{4?��*�K��,��4�a�c�
�]��O�g������+qB�I�F�ÖS�#�?S��d���'�u<��b�*U&	�����ۡAS������ћ�f��e��a�e�H����6��}
�.��^�~]�0�tr>`��`��tx��-�I��T���SCi���']�brR�J���l(�d?}�FV���?=���E��!�{߬�_v\�����B�r��9�o'�>+���XF��ݫ�*�'�~o���B�� :�7�t1߲�BC�X�u?s��~��bn���5?��X��x䘀:���9M�~2<zf�^Ңҭ�� ��o*�^��bU���M��̝,Ԇ~� �3
D*����]W�����
g�,�����
ɭ�%c.�i�Հ�Oߌ/��¥a��>F?�r4ظx����ώ���ʄ�%��Ȧh�ׁ���P�">R}��byL��5�U�卵���s�"�X���|7�-sNR����f_�z�����FI������ys�٢�߽������b� P�X
�G�i�ɔ��M���(��Ń��Mp���f_��c�����~��+<j�ޅZ{c5llu(��R~h��阭���b(�t]���T��7l������W*�2q����rp㦿8�r�l8����1�Pp b�t�@�k!����\,�I 8��3ѓ��~Y %� _�����_.U��ϱExH#�T����XG ɗ&�w��=w����?4�@�mg��{�ŢB�M�r�l%�(�/R�CY�κ7	oMl���0������g1�d����ks�K�0��'�)kpy!e��̐�*װ��^��`���:���{�x�	���3s0?@ʞ��tn}s�Y�<Z�/\P5a9%{C��p@@�Jg�ܙg��`8	��	�h�ƒ΅�K(�4�ު~�aAw�e��@!@�}��^N�Γ\�}	 �&�	S:k�����T�۸�	�<_���5��b&�����W�NJ+j�����b?R�F���t��R�!��GF�a��.�������e�> �ث~���r�%�.ues��#�z]	,�D�`�ÑZ�B��q��Y	jl��r��V5!�7<�7	�V�IZ5-�z֗[R|�ELԿf��
ι4�F�/�,#�7["n����xr�OZ�>ҕ�%�����~
��$�,�2ob��?s�_���IK�A���y	�� ��䲳w���R��	�U�3,6i2^��V��+i;Ұ��O;(��N�v�V0���2�%/����ܮ�BLJ C�RM�ڡ��w��������p!���>ش��|�y*OÖ�M�5�WHt4�ӝ���O=��7����
�$��L�X����s41�5G������t���(��i��}��������46|X�!G
�
�=��%$%T��P\O�i�!��®Q��
<�i�����S�˺qu����}�&�����\�(]��	����-L�]�-�G��6��i�?���ď-V?���'5�R�����)s�����S��x6.[�Q=ρ��o�u����.�Ni���?-ɇ�%���Wi�x]��C$4k�j���Ih����<i�YfӚ(%v���a����r%C�n0���G��Eo@Ɩ�юfp��`U�~��<�f�
�`<��-��SPC��6��?\�fH5�O:ɣ'�Vt+�����I*��b��z��g!�O2�+A�U�S�.)�S��)_�Iә�Y�@�`kLȦ��~K�`CCA��S�dDdyq^��N(����j�z}�ED
�^�H']�!��=�jlX�tׄ�@,�it@�=Q_�@Ev�'x�J{J��&+�Ӯ����M�������b�5�}C�:���$ZQOU��,�8l�j��7��D���n1��p��*�"KjO�=��Y�W�E���nze�U�Q���4~@�6����o��M���]�{h�/Of��.��g_nD7A��Э����8*��,�J
�(Y#` ��o��|T�T�aC��� �$��%Ŧty���n����[�����Ji�ӭ�(�1���@V+�cR�v��o���f�Ј�4iU�0y�	X�,z�Hq|s�f�_)��#�6��ɟXսb������\�<��Q&ǲ�ч=���-J��	ܒ�~��-�6qءh$ɓ��������I"F?���� Tw>�+@|\JvZ&�pS�2!���kn���L�}%P�B�ٕb�?��v	�  ���<�}x�ؤ-�4��)"kOA�V�F�����QIЉ+Kf:?��C�"E�i(���h�0��.?p�W�{b��;�ͪ��y2��O(��V�"hj���ߓ��W�����c���T��kI:BHtDs�y�RsV;ժ���7�/�v����nњ5���<�0D�Q�Fޤ�*;��.�:�,pY]Ѣ��M���/,��,�A���m��O�(Ƴ�w:����{!�_��z���n
�6]�\�+$��^�Yk&��}����R���bETĢ���V�̖M@% ����[S}�ص?�n��z�|�`����dEu�mP �NM�~��i�l6�����4W$��6o�� (>�ލ�ɛS��ϱ�7�;�����!4��(y�o`�nw��Ս�,�2� @%��/ЍD̬����:jɂS�ݣ��7V�3�d��k�VN?��{�Q��4�E:����(��&	&�0t"���e�EV���� �@-���*򾺐����L@29�Oi�yd���K�)�}��HRQ� 2_'%OϨ�.nb&���K�}(w��Rb�k$o7#�D�v@x������L�vē̓�!��`��S~Ϫ�����d �Ln}CV��Y좃�k�y&jL��X�w
ysx�](0N&���l]���b^(�S���T\K�&w�*R�{W�둯Ro;v;�0T��!}����O��k��?\S'�o��i7٪�̣�V欅�C�	���C]�У��N�)W�l�Y�+֓�}��Z�`=�+!���Gl�lt�d�wm�iGP}�*� ��{b�+I|�� E��n��%�Y����U�];� 2�*yH��U�㑓���#8���i����X�%�b:��5LH�� ����F@��X%Oj�G������SR�.��������	|d)Q�D��f����a���$L��&+��Bj���'2!����~}L���߆�)�%!_�a�<�&��2��
��FBr���!����g�D>����i|�p��r��e�˼��H�9v�/������I���cUd1E���%� 1y5�S�$�5�_,*�u�Ȭ�K!�'Jz
��9���^�Ee>����>:��s��`��hNC���Q�ku��6���m��\EܠmL[ ���M��c;��Z������5��ZR��pؿM:�>1%�xNO�������2��0�	`Yfb��@�&�j�rǸ?�̲��sd��<��}���w G�b��~A�¯8;����<R`�~c'�l��p�)��Æ�)
���i=��,�	i���}QjO�l(�������W��Q��KyƸn|0�	���FJ�J�3��_/���J������ v3�h*�ro��tY�g�y�|/>-ո ��F1�p�\"�+U�z�"E�)�5�"�Aق�����,����B��j����{�:��Zo�D!ަ_{L�$0�|0;�V�q�v��R{����]��$4����m�QQ3�
T���&df��2�+��w�?�د��t�K����K�E�ҸtV�747YL�?�'�Y�F�/k��/�L-*��a�A�LX�-��-��32��T}��LD����/῀9���2�x���7����WΌ4�V��׵�X���L��l��~�B��
b���}��zw�|�g_#FV��)gT�[�&��Ŗ�B	�i ���(���ZL]���<x��Q:��8��6���-\Z��&�[7�C���d6��=h�x�PWQ��X���R��n5�_��i���6�5fL�E%ǖh��k��ݾg\��!�YXt�]�d+0>�!��i670�8���`:�o'K��%���fO�&^i�P�]��	a
�K��q|�F��������S�В�����0�f���/!� �I�zT��q"")�:\�mF0(��� �.���!���I8�e��} �# �-�N���IDo%�Ҋ����g�8vZ��H	���F�`՜u�K� �j����Q��F�\Q���)P���Z����a	iCKf"�H�6��@Z�G����K�X�(tEv�?�2"�'>�L��?��_�#걐Uҧ�����jO��!O*Ձ	A=���&]�d��x�KhU�:N�D`&��3\�w?�NL�� k�F5�|?�.6����,���'Jh�dc�H,�
�5����G~�zr�`� a|^JN-=H�)�T��������y�$! �:��� `�2~���bIC�Er֟R���ĕv��<�/m%�`�R,U&����&X��U�7���v���æ6�@�0#V�}�[릎�"Fϵ/�&K�-#���iL"�٘��i��Y|,6|���aQ8�tuZ�*���	N��R���|3��,v���5�c҉����1��C�i�����h_�pC|7�?��KH*P|=7{qM����\[[Ռn��1�tn&��$�����~��t%�2rM�(��ޝ��ZkT%�Q''�y.���164\BB��G�_�n�I��bA!'�$����hTm��\xv��j�,����:dM��{ �4��g�E,�RP����Y�D���bl��- �E�!�f?*QC=,���<>wM�	[-!|4;RB��Ϡ����_��_��ys[��`��w�^��l;e�&#X�҄�٘!��ہ�������9t�?I�n{���6��<����ꢡH��z��}T':pp���e��R���rVӽT�H�8��}�v���]��-Y�̂3�\|�� b�q��\�P�i��6��'1�JA��}��=��	�]"���<�|���Inx:�`�������P ���l��A�zh���9��q�l"�|k�(F ��5áe�-�`7�� �{ےzF5� yh�����ύ�K��?�p�f+���zh-��H���w �֎������g�ݟ�J�i�βG,淆i]������xe�1��^�敜ܫok��{�����$]Y'=Qs�mw���vk�)��CMR�X�܎?y��R5�|�"��Ƃ��$A���Y��2yydn8�5�eIi\~��|9��k�������bJ捨��ИznT�6�<\q5k������%3ƉG�K�*���ޒ����>��_�|Z}����l��Y#S�e#B#3��8�``�t�vd�avB%�#`��~���M�B�rt�$Tc���x*���1w�4��)��j��,���O������O���_�$�&o-r�'៨UZ"�5��!̵�&Fچ�o"���/��ᾀw[��u�;�����:��p,�(}��/ >Lg�|'EW�f��L��܊�'�2�>�k�kϦt�UD!x��.&~�ݰ�u8;�~[�L�2��	�^���Ry����s��H�s7R��������"|
aݚ������*������������4���J0A�Xڨ.�"_8��f�^��3@h�9=�*Mf!�9���
U�&����4l-d�H5C>��B7�C�54�s��x,�u�e�+ZơE%���z�{a٥��%���r(��۰�dLն=�5O�/˔�Cؒ�PwB
���~���w�m��y�񦸛B���@ն%�
�����M�`}\q�=�u�����`˅c�����.���Hu
da쿤��g��]R�A��v�L V8��kف�y�P��Z�bY��B0w݊�4�9���o�������W���?�*�kK��h���z�y,=���.�����QF�>���}9'�-פ���mH>R%��j�jTKҕ�e�)��$��[����[L1r@W������@J	��bV�g@_��'b���e�-���� �ݱK�.p;N��UHM��Սn%��#:��O1S�[�"�Jd�߆F̓�3���S�P*�"�n��;������i۲�v[M�]�Y�nl�0����۩p�Gv*������a��EY�׊՝d��Yi��}t-h��^\��)�ta��E?��(*4g����ާ����7�i.\��a�o@����n5a-�XXag�[C����~��J���+^�u�L�b1��ɩ?Z�L���fB#��|��إ= ��Y����M���)N�٤�dp��%�z.!Ý�o[]­����m��Èd��s-������z*y��M�8p��a�oG����� ι��ǌ�Z���a(�]�$�6JNˮ�� �ح��
�����u�T�By�c��*�yF�B�:i�%�&z���}��S{Wm�j��p{��`bM'��c��Ó@:���#�D9�}ŨL^1�v��@��v�UQTq5B]�R�1mNʆ��,��ab>$��,h����8u::?�)V�ع�����P^i�->��cG�I7Gv���Q�$����<���2�%r��F�ԅZPGl>D�,SUP&}p	�����|����խ���*�r�F~vWܭ��!�����i���j��4X�Eol0�5�J��N1γ��b�x#�����GR�VR7U�5��3E�?i�,d�K��Rme�¢3�����C�lv��M�/��R	����׶q~궏{��,{}:��`�揜>�ɱ�B�+�.��|�)kS9�>}yp+�y�p'���vD�Ħ�f��m]�wzOa��ȉ���L��*��dӇ���D&��B �X���H��az#��F�c�:��=���x�ÁU&�O3�(��'KV@r��o���|0���N�!����n.��8Y�1���шV'�\q
����jb�8��a�7��1t��$q���/��S�1�=�����~��>VoY���`t�ӗ�79E�J����bS�����g�:�->#�e=_�
��Ψ����/��?$G�QkNJ��aL��1�m�}�-�����'lȐ�z�Tq;��WHϞ<�5B@�Eҙ����N>a��
E؎�Q��h�䰈���I_����,\`��hۅ��8����I� �:�G.>�z�_�aѯC��s�x4)��Э��8�ȥ(<y��A���u���j�WӔl��#�a �RH��za���*��.�!"f[�ܓ��6����/�Vm�.a��Yr��-6J��:
�KI:�^(/�v�l��+-�	��}�Y��z � ^��]�+b'��++��Y�e���\�2:��(���'�����_Ut�~B����&M��[�m�&��s���nb�x���0z]K��1�Vl�ek�`H�S��#�#[Ȗ���^(��~�I�b�SQ�,(rȒ	���@��	z���L��('ȅ�|E(�$^��JYvR"���
y�a��9�>��n�I�.�9� f�P/')'���w��	��ݲ����汇��~Ŕ,��M���>����g2�K�gFH����5���6�k�P tǈ����m:d"~�*��د� ���F�႗{��=2�0����@)�i?�1>��k�̫z'8%�3� ������{��l3�>%oW���t������D�b!��b��#�f�%��b,/0 i�ܪ����=ֳ6ȇw�bh�������^aV�$"�V��4�`������2���d��p�j�p�+޻g��鑔�VEŞ�DMg��E�]�2@)�)���7;P��D���5���;��,	�9�@2T�1T5�x��<d�Z�82��5
N7*��c�F�s��k��6����*~�"^f�p�T�/��{�FR�i��"b�V|���°Ex�v�}^[��]�
�3�l ���̱Z�������w�����YM��k���nX����3�;���ަӂ�@\�U� ?v�+������J���^na���NZU���)�GY��:Y����JZiJ<u��p�bUC��ѳ�.g���(t<rs�&ܵ����I�
~�K�t�.�����W8����'�$��"��ގ�qȌ$���!W�ߑ�ý#m7dC�(�������P��X�SD:�� ̊d03r~�������� ��8�\��1���m���ݯ�,4�<�����������h�r0���(V���xI���!��rY��h҇ ��� !�ª��C+�0�~�?����l�a)Q�Q�=F��ײ�