��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%��c��g�t嘘o���Y��
~��>�2x� h|�tup�Xwx[�3WD3y��]�����Rhm�t��f���p��@ށ}%Y��j`r�<�{��8��LN>_��� �݇��r��U89��@3�\	�u�B�9f]:n
2�_�1EL	�K�����-��i��Uf�K?����T��f)6}zFŹ��@���ftt��{���u� $#_꠪�iu�aS�cm��a+�m�e�|�J꘣CS���l����o@�#��w��e����;�f��]��Xoa4柭|����_t�=w��A%q����it?�S�t=���c�$&t������י�D�@�J�/��(e�GhKA��W����|������e������q˝В�t+B�}wrzx8������n���Ja����g�����NmK�d$�5\��.*b�ǲ��7-i&���E%�VΒ[�)�����$)�u}E�z���=�F6���?@��+������R����{FG�������}�*qU����>����]�b&�s�R^��މgu��<A*��v����������D���M���F�ށj�|�#�
  ���}0���ӯq���ʡ���h[�})��A�}K�٪C�hA:4�Isr� ��(fV�_�F�z\�Q;���@`��!s��{�醇��x77f�K��E�����f��h��P��H�a�� �D�����W�wG����!�-a�ָ%b��U�P���t<UFa������gj\%�$������g�Am̿-���u-��2ٙڒ���I�����	f����ٓƻ;��&^�CU��_ED!�k�q����o��u|�2�H^�S�n�!��C�4��&��RVJ�O)xp��2 �ɥ|�s3×9�S�*��E�.�>�_"��_�T��/e���N�gڶ��������}k��C&_&����L��΄ �מd��x|�E��F�tM��R*�+{j�`R�F��7Ϭ2o������P��u��>r~��A���?��=gG�P�� ���}�΁�U�]����J�p���F�-�j�ʻ8�>�i�li��͖��'�� ]c���h�G�J��K��Z0�SxHb�"A�g]�
EU��8t��&2��O����$W�s���i)�'x�J
ST+�Ѐ���$���]VZ�A��~�z%�u4$'��28��KúB�+�zX���m��·���~�T�f.E�T���:��r���� ���t�>�R�
iX3�^�r16��vf�ᩄ/i�	�▞,'��ݕ�~�+�9�Pm,6W�����q�\M�h%1�o�*��]C+ц(a�OG���:�"��y1�l,<�Jgsjh�Ŗ9o��I�C/��*C&�VDj��a�fi�����jV��R��z�*�[����un��kz�?���Ujc89�䀐�>Zc���殆�Ci�Bm˝��@<B������6QA)�Β5���9��Q���hU �l�{!Vm}M'�!�~�Nu�Mzo"h=4��h�xQ>%w�c� �׿�����E�����W�1��A��� 咖�@IժXEz���7+�ʇ��?^P��
!��������/~R�+Vj����˺q��v9j�0�=@O?���*�*S�,*�!gv!/ե��,!9rڢ���d��]�Y�u  O�TH��"K�Ψ��Ǵ���};LC'�0��B�o�X��<��ҩba��~VI�� ���컂ΊU0��/�h����*/�?��p��x y�ӊLo`n�������/")u�Y#���>���z��*YY��b��х���k]��<ܖ���-Q�����2��������fʼsL��n1�Z��l%�Y߂��R���{I��z]�,�20�!��C@��H��رʎU��d�-r���������Q�:������VZ�Ɯ`�"�������J�Qב��=�U����v����\�����5.����{%r�أ����1ha���b:Cw���X�?����t]w�8&{��D�I(r!fX���*e��Z!HO���;��h~ѹ�)���3�����-/J����~�B*�)��;Q���%4_F�CK�.-�Xw���a7�۰��pB+�k,�c��x���a��=�;��\O������������❎�	Lj�v1bHH���U���t�H��iUp&�E�g?��+��ϰ814����o~2	�4��B�~˪���YʊrYMEl��'ז��v��s�쎯�莱�����'��E�P����ɫD��Z�$��aO{Z6hîwP�a($*l�����"����
E�~�{$��]�<�;ަ�
Gq�˘��F`��uOY)n�\Rf�|��.Э~��ԗӧ��1֞n�cj�$'gblCJ��?��g$�/@���!��IR�ϾCD�����:y���Bݣ�GnKc�ҟi8r�)���6tO�!JO�9l��(���ʪ��;9"�.�q��Ԭ�ٹ=�.����#(�{�J�k�ģw�xH�c	�G�M�y����(B�Bh�QC,���v�y,Jq�!l�p�ۼ�iԜ+��b