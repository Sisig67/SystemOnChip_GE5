��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_��՛	�D
�T�da�]L7��~yR�����*̮AņK��+�3>��0�SL����.7�S�^�E*�>k����l'_et��f�5�����e�t�cց�/�\Y1�>=G�$�#�=���7�B2�O�Lb���CMy��$n�K4��iF7;3��j����abX�t�}<Wy����:`��6:���D��%#arq%�w���B��mf&(�j.����F�vZ����������	u����8��X��J�T�J��P	�6��xD���u* �O�S�K�@_(�sX����zx.(9���E��x@��a���Mdv�	�q�s�r�'� ԅg�a��6 i)�����P��0�_K�B���T�k���c�Z�:��2Ԩ�A�ND�������/"Χ�s"����SP��jN�!����b6>k�nWXe�eϠK*�ɼ��ޡ��Sm��)��2�aQ�B8l�����p�7����)�O�|;�I��V�T=[�&�<�k���5��2�[*��3ҋ4X��@���/BȌ�Dիҭ���Đr�zS	���uH�}�ߔ��1~F���"Mb����#\��#�mw%�ƻ�;)�y��_�̿M�pmZ����8&��li"���rSf�Z��X�iTM��ݺ0��?�d� �F����9H/x��|sm��6�FBz��xV?<��������ܻ/��+"��.���a^'�(�y�ʷ)�y�S��.��֕�mo�_eU�r�mk����)��e����9K�Hϫt��mgoeMB�g�� �HD뺏����!9��E�$�֊�#���b�u?���qT�ߖc˂G��u{H�|�>fd�t��Wܖ_�A���xQp�
�+�2�4κ+!���v�t֜&�ؾ��Z]�Џ#��֋���swm�(��P[�֢���:�z�v:�CW�`�r>h
���]<��ি�/]Y��D�o�c"��4��qVAwf�
�<� ���I��C&ͨ�!�2t��(����Y�U��٭��h�y��4��8Mt$�Z۶ʭj-�;T��*LʍV���^��,�B�:J("7�ݗ���D/�4"l��g�J�Y'C�gp��ct=J�����y�W�����H�%	[��VQ�  Gc���Ewn����
dȌWz��ය�F�Y`�%�=V�+ެ�h�e�G������3��;�Vźg��|�C�K)� _]8=��)e[r�U���S�<f�X�,7��}_7�w&���%�FnQ���j�Aw5T x�S�����49�	�{=aeӕ®�?�F���0��ݵ�}꓿x4&�u��
x��V��ɰA�i3DmM�Xwi7�s����!m�P�uk|���4ew=��.���9s�_��o��eO��R��Ʒ�M�3���Po1ZR����/��.%�R���X8�#s�4ե�Nm�Eh�g��F*�R'uG8;���x8�Yއ�;�l,nܥ��;m$1�)��E�W5||@:�5m�/D�F(����/-��"�$\��H�|�~D6ȑ�_����@)w����Q�m\x�M�@�U*��	h'N�c��_%�/�PU��9%�5H����h�����X\�<�S���$��V	�Ϟ�H���x`k�d�͔)���a�����[��Ş̋y��ѵ���������u=�o+��ɂW��/�O'@g�B�Ӄ��uo�� P�;�H[  #Ŀ��G�^#XI�J���P�\_Ƙs��@�;����������V��y\"�
j�.?Ph��<�gE��dt-Cp��:l)p�	��E˅���L�|��xx: 	s�������+��������QcL�<ե��zVJj�;�ߟ"�����,���hk�W3���ۄ��52:�!?��U�s{���1�OO�,�h�	�0�ztLoĂ@�_ֹ�I���6O0/�G�ؾ��a�����t���ּI��(a���J�2g�0�r�!�]Z��{�&��g_���za���Þyie3b�1��F)R�pJG���o,���tW��%�CJh�4�y����xyG�_��-N|���Ŧ� ��ʃE�#�[rQ]y�x�,��dm6���-/[���ǂ��u�CG��F������m�!� �]���fL��B�$�5r:V?�r���ay�n���o�.{�-�mkBf�@Y}�|��](&�VO�oZA�>���':51[	I͏���\{�v1���;��v����/x��"��O��E^^\�S��q�Z���vM��*#6ӽ�7��2rw���d+�N4;�%��k���62EpEݒ?l���A����[V/��j`99��B槵?��x��{��f�,,�
���e�	���['�3�碈[a��H���\d�&�