��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2ic6�Y�FԜ��m�V�FҲ5�X_<��V�a��L���y.ޑO�О�����đ��e/qz���KoE�`s�4�K��_����F�{��t��~fT��2��h_Î ����a���9�L
�Eqf�xs�Ӈ�|�J��*�*s���n��,q3e�'����-(f��lV�S�R�>�Eױ͗�/O��=GI̚�*f�6L`��b,xLqé�,�_�5���d�u�G��� {���9��<)���tR�x�=�������\o��G��w�y��p�.�tAB�k@|���:�G˾�?�b�b6��
ށ蚿��Q���:�"@���RpϹ<T�F�	d���EA��ѨmT�R{�Pk����4.��Ħ ���5��-,Eɏ��q~;�)$��w?�OE���e�R�Oi�Dg�Ņ�0�Yr<��T�ElKvKyE#`u3�p'"�	���k���9�"x|Z��ɼ�e�����٤!��s�94{L=ܧ^4��t-�~�৆SY�oxy�頎o����:���Ё�C��l����\�5�Ǫt�<�F��qbv��u]���I9<;�����v��|b[U�2��69�Ԙ9\c�����Q���)�%D�5
k��yҬd��.DX���z>��>6}i5��N�|A^F�X6�ɳ�}ݫg�� oE))CYG�X�;Ĺ]:���উSڋ��	��o��hpf��[��q�/l1G�y�k(�]B,B.�I��>]ʻ��0���q6i���b��r_1��7� �>'ţ̨fyM`�k��+i�~�c�R�^t/=�X�@'�j�xS���"j�A��b�g��SQ�RU�F0�j�t�^ܐ������c:��S,�2�,{�;�`a�|��x}/j�:�q�4��E���F�G����h����*CѰ�L��FM�䲂$Ȃ�p 7!be2v�p� ߇�� q4g=�/H*/	��S���g6�x5uz꽒ۆIa$�p93�ˤp�^Gb1P�B��z��	��jj�A��I�7�H��
�t�Uy�ǚ�0��*$��S�ћ����`j лzq��<�-i|s���j4�0�Ʈَ���-	��{|,���xe8,-�M�C`&`�V���f/����ף�k�|nF��6v�#T%`�ª��^��HE�7�k��w��V�i��i�닙���a���9�l�l{�$�l���>*�v��_/Bh�NH��'Q��2����� $�#5rM�J:z�o���Jti�+Y����Į��"��O�@*�ԤR�����{���`�Q��ڊ�I�b�2�J����Ol�q�'+{A����~�>�Ԁ�c���天�J��<x�H՛C��/z�F�(��^�e����!E��=G�xP�4��fCDڴdi�NC��:�����Du�t�y�R#f�qBv~.ږO��)5����X�9<yK%!�B��[����-j��TL�$5��� ��پ�l�n�Y�1A����	$��������5eʱ��Gڱ�ϡ��' ���?��9��L>R���Ij�	C�X��G'�o�	B����D�q��)[k��%m�'�����%�{�z+z��<&����,:;j�Ǧ�UCk_eS�;��F&�+,���4ոR�z�����0M]�̈�?�7��Ȍ�v�қ6�J���]BL��V<��#�_٠�8�H�7l�D�1Ө-×���B��6��1!���*�.����1���G�L��L����3���K̼4^�6zH��&Ӗ�bլ�r�$Q&���W���zK�ڽ��XZp�Ō����^��Fm��2p+�7�Gk��zM6��5���湷zS�F��]���\I�~	Frh~�m�x'n�� ��}��%��Y���T;;�M�J�S���s�3��<��k}aD.7�c��]�m�1�C������f,&���o�x���e;(���#@R�!��G�v��\�p��{���� b�JS�ۢ��0�� /�g��]6iU��[f^Y��w����H dE��Z�k��������6�"x%��][���[藋�HUvzF�D\�@ϛ�gxdڈ�8y/�JH����𓍺_��ٞ���:�MA�D6*jF����8Y�-<��G��9%Ϡ�V�24d��p)�h�/����8�U��V�����G�5kip�/~���>uS����3�Es7�ۮ�O��v$�JfE�s1��ؒe��.�_����Y2�����gU�0Vϊ����D2TN��/Y&O�U��=ٗ�A;pr��ihD�4��n�j�ib��F/���-2�ɗD*U��)ާ#��p�.�94�*�U�-*A9U��ۚ�p�q�/��T|��ާO�	�?���=�$��R��:�*�AK:Y����\���V�
 z���4s��ƊW�H����ި���×��uV�:�O�Q�E,	ozm�2� [�sჳY8��h���ҬJ���׽9_>}�"I�J�����hF	dF�,4 ֥<�g�=��t_f@:R�]�>��qڭ�~�ߢov� ?��	�kf�T̥�d]�BO����:&y����L�_�������Ni=�W��.YF�M$��W�x��£���m��J�
��a^�u��)��\�6��+`ؿ��3�0W��[$F(vAj�u5YYGv�u!�����-X�����������  ɼ��nk�[�C����]y.(ȩ��∾�0t���\�ז�l<�-r��h囖�:	��ޥêr�P�M!��>�)��w*8���}��}�̰��^�w�Y刲4��O@"���|���is��Uw.�P��S����(,!���y�ѥ�2y�:)�ӛ����4@;K`G�Ne������!��ss���yD�щ���ͥ��H��c*�V7KH�텵/��ӈ�+�a��M��-�1����\�z��/ď�t�H�	�^iG�%��-�i&k�n�d��1���H�s��H����f�5�p���_����ZK8��a���g��U'3���L��]L�I� >t=��y�U�X�6r�O�/ԫ�>��|fo.<o�������k3 X1U�'7�}��)�c��p: ����aw6 >�s�y�d��1�
:~O�e�����!b<�i��Gr�*)V6�V��9&��/
V~7��w��jM*[�7R2w��5�O�o�,ʡR�^[[��)U>E(�"�����ĵY}�8*�.T�&1��+�؁-�����u��zIbHQ��kCG��-����9i�;�����qWmo`#�ɽU��b1��K���v��?�5���
�8�z�G`΁m2��>�Ve\�	�V�Ƣ��P%��ywJ
�57	xōF�Tmu0�$I�DqM��oXՁ����;5}W}l���zK.�U	�ߌqZ���Ӷ^#I�t�
7{Ͻ���,,OFתs�Zϲ<�b�T7�:f.�?u�S͏�̡;;�"�n���������R�'�Q]�	R�\�;i6t{��.�!xPM��))��~1��6q�7(1���K41F�n��G�oG��aB��)��m�����E�r��w�;R��(V�F�"h�)���c=t�ܸ�pVL[��\��|��}4�b�q�>������"vq8;��T�#M�,$I//s�p��]<y"]��Z�}w���P"�N��#���9�!�"���3N�X5�;̞K�X~A��N�~ڗɞp�yؠ�R�3� ,{����� �Rkr�A7s[B�ߴ\����*aN�.���¿kj �־w~A����;��rI�c����=��{`d��7�A�_GY���olhS��	���`�Y�G��J���h!E����ҁ�>U]��B'ϝ#���N�f�G��v,򳶗
e����ן���c��6yO��!&��hQ3�	�q�$TѤ�d �SM �`~	s����p3G���(�Ь�̙�G$���)��Q���X�7�"�>�rǴ��a�F֝��oT�l#��yU��p#9:��&���'�ƅjH��gqD�~S�`v���~��hdh����^���M��bΛ^#OV��f�`)4��kx�����B/��=P��aP~ܚ\(����o�:��O�T"ߘo�[b�_d[����8���V`7c�a����}^`����=�F�O�]�H��X2��ܻ�\aO�-f��>�y|���O6��, yE���y	��'KD�\����x�=DDA`G���L8�装e��!3%%�Y��jd���5IY)���p:��]"�۩ҁ���z�f�&� i��nΟ��eʻ��&��P�w�KTFr͢S�C����O��Wp����_7�D�S�j��h)�4��l���VJj�VP�������k��"B����5���]J��G��{�W�d=[�c)�K�$s�m�&�x�Y�O8Ь�F��vG��݄�BBD#1.C~�*�ρz��_�/�@!Qh~��(���n3e�bO�bՈG�)o�~���Q�0�7��/�MX����� ���yc���'!d�Wx��JuX�%;�?�R[zm�3b�ե�k��%S��>	gى��E��Ʀ}������R�GTᙬ��J��������;���y؜*��T�������e���j���wzZZ~��&ܮ�����mG^���6��7=��;��&J��[@��T���.�p��\��4�+k�0;�~�Gw^!���fc�:Ƶ��x-g�1��vh2m�}��
E�:��^��[�ib]���(�)��,�$o��R�z�Pe�,�:I]I�s��)5�R����\'L���c��BGR��
>cB,�h܅�/���{�n�� ���o�sCɆ��?�58����}���?�������^���w4����qFax]z���a+5�l�ũ�F�Ja�jU-B.�w�n�O[��.]h��Q�f4�#��Z�3��*����_�%G>�,9����Q:��۱�'j��{��CR�7:ɰ�]ɐN䱱^>A7�1W,nc�ߢ.՜�,��/����N6�������N()-Y;p�t���5e�9����?hnΙDɀ�R�
>WV�`)f춢�Wb����Q�zo�K�)������QZg7�
҂%(ǁ6�9

���̤���]HK����o�3�����:�ʄP��oJ��|���\��Ƶ2���� �����Z��d谈X����<1R�����<Z�1���������"�6��4��gU'��9�<�
��2M,�3���qC"G��Tj%�$���}%�;��#3G��UU1�晵�K����2�QhiK�cx\�ts��x ��� wA�2�-��B�J��zM����3�!����+�v�U�7r�Ŕ��6�+F�q���0%dqK#_� 6�!���7�����0)B���3gt��N�6�g%�'��9>���j
-�R�B���h�i�<��¢�Q�l=�h}믗�L��i��G���Wq�)SI��\a �gD�T��-���X����;m�k}�e�s����9�S�1��j���h�J>Oࠦ���d���E��uv�ɻ)��iu_m�y#U�ݍ�IGh@^Im`�9С���;e�2�0F���l0rBwQ���fgEq�C��.4\b�Gq���3�@@�@�IK}�{b��$-i1�qb�5l�<$SVusfY�_媔���u�L�����m�����iD��R�a�Q׫,�����P%�eKϵ�10��{�~����{�c�_O�m�Pwv��q�>���/��!ƛQt�����6lk��j�� �/�T�'g��瀥�nZp�=N�PD�XT�ѩ��3yL~��Ĝ9���OV�������������D$?6օd,&a	�g�:����Q� �� 	��72�������}�w*�tZI�kT��?�^k_�����ޜ���w�������B3�=�[���������H�i	��#��MdK�Z:C�+;Hv���K�^��� �;!w�ߙd�CTHѵ8
2j��[��*ӛ�]xYmzG�Ҷ�NW�<�X��#Y5:�g�bڲ�%h�_�x�rc]�p��({��� F Z|c�,"��D>���P�B�'���0����X ���Y ��1+޵��DlT����c��Vdɒ�1���~<�cӈP
E��C��b�QKh9s0�Zt�['`$2�>[zna�Ǟ�$z�PK��"ۺ�����PR��*��{Jtu1Wh��S�M��m��ƺ%�u�.[����ސ�}8���r�yf��	�k�M�Y��ˬ��!�0�O%���i������$�$A����84�be��@��%��� �輞GR�=K�x�����M� +p�H�&-�>��u#���׬�Pb�zj�`\�!��c�!Îz]$��o@d��^�{�|7ʒO����O�*�)���}��;�<��;�z`�3��� �	^�B��w�99� h�h#�ۨ����a��S�\iAU{����7 V����
���r�'l�ͫ��_�^�k�n�m� �Et/��	�6{���)���-K
����p��8s%�1*�3�#K�D
wt��IR?�,[C��%��n�gY��@�ͩZ�E�x���g[��gP���ٞ�'8!.1c���ƗrRt�Bİ� ��j���u�7�PJ����`0�Ur�a]��o��~�@�4�pj��4�hܴH�p��W��SgX{~w_�ߺ��t�[^f׈e^"6���1rp�<��P�N�W���?�܋:j�̣�l
8{��٠��Іyuum�{�}䪛	,���u0ow��ܡ�<~��
��l6yK��D8lA?�������h����'��/`��N��!�M�'9)�9����Kwݛz�[$�G��̂X��&]Xx�e��N�����Ƃ��UO�Ȟ�x�ӧ8�Fk��LЀI�ⷭ�?�#���Oy��!�����@��1
kbcŀ�ZG�ώԷ�>�sY/T��u����\1�L �ߢ}��Z�>X�:�q�k�d�>^ZGf�/\��o=�$��P2���	�:.�ߕ)[�b΄��3 \w�ڹ�m�Es���Vv�Fu��(K��/�JN������M�f2�'�
7_I����%Qb�oT�L-tK�V��֦4��� <���xN���m?n	�h����q��=zB2͟�4褿���Q��?�x�3FS];I���g�o�GI�\j6�)M��N��TO6�7@V��s��@��~�����#6�k4�0��R�"h���j�Q��] ��x�p�`�.0�_�=����QԵ�TM�P�û�:Vi������t/@�|�������,��U��
������޳5�����4�<Djb��A��.�c�K��2�\}}(w����U��ܺ��y(Y�����Q�5]�>L(�/�+6�S�S�"��j�Tp?�oU�n�K��.�uA �6��o��G~�D��[IfG����c��)�ߘod��b�7���κ�#�.���3D��Y=��Qp��&Mշ���4�������_��
ybm��d���v@O^6�7��jx��?:G\��?�U�k�g�@�n�����j�̱��/>�yǡ�W�R+�q\����o@a�<�V�@�	Ax8��ڸĪ��P*�����`���g�����`P�VT�x�Ѭ�� ^�YY�1�>}�g4d!��s�C��\p���R�,����h�+ɪ~���\��*&/Pu�6,,w�3��|-�]|m��փ����Q�4H����<��^Ǯ3��e���m*h�Q}:6Y؄�%��,A^Ѯ	
=��뺫�lH_0ǲ�G4��0��I�	z�59H�VO<?�8� 8��g\�?���i��?DA��o>.H�������,y�wl|��J�Ś�i����F��h'Th0�F�0W�|��<8s@�yM��k�	տpk�v�,��0����:�����V%1CQ�>�q���VÏ2���5B�Dz�Ӳꠋ��(#��V�;��D�{(���Eڜ6⛷�K��(E	�_H1���'�-���o�Nx�T�РW=��hi<�3��54��a����CL4s� ��������&A�� s�"��H�ߩg�� ���������E�u�ǜ�Q19'}q�����v�*�5�H �@_�J��4��t�{�L�7�^��m[NAE��ܧ'�C[(Ot���C(�g3`O4������ 8SC
X9%6�ܜn�8�#x��	!��	Ы�1��$�N�� �1����YuCS?0��(�:I��X��D૤v�R��,و�p:�(��O�Ѱ��ND ��	 ���O<O�� vX"������
�P�%�*�̬�����u��B�Ζj���%낧V��a�-�ƾ�x.�{Uqs��,���
��U+��y �)͇hf�9L�骊�Zq��#��,G�f.�q>
0��%�����2�)%P�K�7H]� �nW�	��D�� �`G��Qj���&�@*� �&�V���z�^���<��1��&�Tѕ�ퟲ�^�w-�"�������=���9v�]F��$��t���ݹ�������@�vh�I7��Z����FՈ���y�7�bޔ���n@�I�=m5�{B3̅R��<E��F�����8��4չ �Ga$0�&4�������c#��_�1���:�)��3���O�hwb����$	9[��x����	����Ղ�c#�5sZ^��Dj,���Q��~�>�8b��C�؍-��pZ���H�$TQ�t�Q��;�@�N5E�|�������I})h=a�"8t'Ym	i�?�q3��"�Y�B���]3���I�70A>ZT!Q�I�Mk���c�u��/̺��K\_�&�Tq��P�qU�hp���w�לBw��Yy����>v~��Q] �C��� ��>�<n�É�q�s�ܣ2�X��%�^F�ƃ/`uX�=����$���*���/����l�ńa&������_H��g<vA����ob5�{��ֳ �B��j�J�>���al	��*a�P��I&��NPsw�J��
$$y����^~�I�!���CR`��R�Q���m�f�	f\�Џ�~�~݌v�:R�Qo����o;3<�p���:t�'�@����Q���+j��9��)R�rn�U�����_����/м�Ybh�;�f|��Ċ�{^<oQP�z����Z��������q43���� �q9w]Oge�q��8v�P�o*��8�o���_��[�`G��(&����B�㏓�5�C�3��Y��l8����n۞��wk:5�P���TI���H)���r�"���~�Ԋ�D��O����~�+^Nu�r�څ$v�� W����>YSK��.IaY��]#�>r
ٛ��~�%�����B0�H艄�o�S����a��������ݥ���9GkB�ic�u*꒎֦���d�o!Ŷ��Q���޴���⏏��6u�2B�	<���|���i��C�V�T�/P�|%��\�:�\�:\��Fy���B�5�x���{�{���Bx��Q��	m?�2��Gvö�c�&1�?B���5H��ni���	3+vZ��3E.��꘶fZp�|aS7�~$���)}C_34Q@my��E����m�ȋ�XbeF�
+�ı�Bܗ��k�'㌍�>;�<DҰ�<:N�F��yV�lM�k �߼�LdL��K�9�!�n��,6}ꖱ�������O"�cC���I-9���I�hð��TѾ\���d���C��o��^I�ET�/Y�Z�hP��6>����H��jPp��>l���5����Z�F�h�:��8�tH�Ϻ�h�*�9~�+�D���p��I�!��t���H��І���剌=��ɺu�6 ��(��I ���`#�0�3�M��0���%`�d�0�<G�kk9x�7�������p�g:��(��Dhʷ�sdC�Fl�ZNC/�/�Y[��x����b5��r�։�9�E/� 8x=�m�ݬ� �v%N�f�B	�����H�i�P�2,
��e&��C�=	����0�:�I<!�pT�!�M&��$�_rvs����Ҭ�{�h�|S��N�Z�6+9� ��U��hr�Zcvy�t7�B�pq�hݣھ�Jl�h���u'�7���m^
9�c�4(>�R6$4;�6�e�,�M;��9�����G��e�E���_%���	�@b��X90SV����c�� �$�8o���P��C*�����5G�m���Q��;�ϣ���QL�`!��e7ZFE���Y7�1� z�K�A'�]���u�W#�f_ǀ�0,��YID�`��f���C������BK�q�+�+��d^�xS�{D�ReuA웁�%j�BW�\p|������P/���HJ|�(�0�A)�������L���jǫT���)W�&���\��W5RH�U���� s<d��=�n���ip�0�j�%�X���r/�E����T46eg�d����n�����Ï���>���5F]�RPKP1�*��Ư�=�����~b��p��!#��rˌ#�PDw �Y���r�����M8�>Y�pQE��!7_5-@ �'�9fզVy�ȭ��	�a���{��竁�4:�����)��L��!�8��
�-yW���l�1�qd����,+n�~��V��Y��(����*buh�'�+r�vz��6�T˚.���m��MF*��{6AW��T#3{)��/�(�fN�9w���0���H�
�4�_sUQ�-�8oXF�̸�x�ճ�oS�6�׏�u�T���."uyJ|&�E�Ջm���-Qșc1�ٯ]j������6������p3�P����8���ĐU]B��u��;�����H��}c��h�K	�����J4�j�#�������_տ���Ha�f�'r�s�T0��R[�Iv�����:�Д�E��a�d�D4�9��
}���A���9�p�{9��Z8ڡݶ�`	�5e� +����M�"H�][��� iD��@G��4�X+N�%��n�e��I���먆�U�H���mv�bmA�f��gXF��B�ʎ�M=���`ԞvC��9�1����X� r@�%5o��lxN��h!�F���v2j,�E�+=���m�AFs��$Y_�q���`W�;� ��#�]�����#��W���,[�,�;F���:���`��c�vӮl� mf� �(���2�W_3W2����jdPr�3�8X��7���Z��t�q���v���a)j܇��HcD�����q:H~�=�����hl�}��B��O�N�0�Fn�s�`)D��;*��D�C��u{��"i%��L!�&ߡױF��H�-��5���\���^ᯤ6��>c�ю���x�܊]:�b�~7�n�[�d�пa<S�|����I�iNi�Ը�G��G2y��B����`u�g~�y �z�~�0����3�K��{�^U�Յ^��gApL*�������8@E>��B8�y�TN�Xg)	<Ҁ�vT����j��UWN�Epp���*{ 0�ªh<�O!<���5���e3D|�8�Z�g7�Ř���H��.t���?��[L�L���'ㄓ�����P��y=GK�`�s�<������g*qO��o�ږ���hӯ�t�`9��G����P��p��ez����݃b��iU�yF8��,p=�D�g�2܎oQQ�r���)u�����p���}¯tb����> �@�A�Y%Hđ=�v	_�z����"��]��څ�=`�775����: �EIa�Ik�z-ݥ�M�.�N�:���c�藈�|q�]Lka�E	��?jzZX�-�H���xU��1Ɓa�]��b����a	�jV[���(�@�yk�����%�&����i&��K�gN��6��ʊӞ((V�=O�>�@�E'j�#�e�'�ą�1�OAb)c�� <� ��5�Č��	�~��GBf�Zni�`�E=�H���!If{ƕ�bK�@ϡ
����d|��G� ��w9:�P���m®��ߡW|�mǇ[��Z�F;ͼ"�U��+�}�q�!.����(�����R��V�p�KT�ʹ��d͚�M�VD]ʉ�76}9��YG�	q��)1���|�8Z���A��v� w<��}����{��� �|N��o�5<D�[�L��'Mm��,�
{��Q�b絗���o���G�����><��F��)�-
x�?�d̝"����K���7TA�#�%�ӧqjM����PN���#���j�3�}d� '.E�~x8̐�lq�����L&�&M�ʧPu�`��K���:<��<��Z܌����f�A�R'��F�:D2������㪦�3X�]��5�$�2K�T�����kŸ�Ց�+c ��R=�֤/�&�h�D婛��R#uI�#��F�8 �����2�)�Z���ij���:<�����!�L
D�$^M���ho �W@�Pu�2X/(I�1$B1��j�^��(jyvց�<�$��CCEk��I���@)H�a�����s�"��5$�r�W�Q�BX	��=��*����m�~s�4<b��Xx��1bgu���CGy[��C�}d���]j�ɵ�~��Pǯ��K����$^
��Vع1k���#j<t�F���A����\df����y��mN����GO��Z9c'����hA��R��"A:w..��{_��s)�9`:V	<o��9�ƣ��+�����I�i0&�6�ӳ��(8�DMN��>i�?����]p֋ŵ��i�CR7Lv���ߌ�%+2|rɷjN%�s F!��E���a�<eXe�8p;Ύƭr��L����+�e$��;�@�9����QZ��t̑ߋ$U�&b�P;�'����f=U]��˲�r���ny��R ꀯ3!@�`l�?����Β���S|vzO�8[���殯�μ�;产�C���<��6�Q���������ij����@V�����SRh�+��Nؙ�'���w���C�U����5p`]^\:k\��uK<�i-$�����`��Y��[�!K9�2[%�0L4,2C��tm�9�}2�+=`I�����g�>�n�_��ap:f��	䫝A5<|�f[E��+N6D�K���.������7��jڇzSPQ���Ҩҗ�?sF�,?�&������2Wǝ�}c �K����Y�}�'SVx���!"Q�y�H?/�/�2�Nh�,�������i))�����J��0�l۔�Y�r�j�ϥ���Z�5�2��y�nY<��H����p�u^�d����:
ӯ��� a�*�:�o�v�~ME�_���
X!UZ�����m����N�Gk����n�w���'�|+�+��`[����xH�Ѵ���[�o�^�_X��O1�|�;|�`Ad��Ѣ����W�#d�������Ȱ��� ko�`7^C����k�C�{�����c��uQ�@�Y{n�|����k<�a?�;J�Đ�Ra%Z����y %��xs�� �뀳��S��j�މm�+��Ch��᷇僩���I3�XEa8�vhN|����B�Wrw�aK#���ln�������|�E`�i�������%�}�<Q��#b���l��~��٧�I4rQ4�E4��Y[����4�� ��Ie'�%���X��l�� �~Eԃ�!�Wl}"b���:уY{# c�=�&���A*f=���|!>@1Ck�+�k�]�@d��T���w^v߸ИY�#G�y���a�kB<דYT<byBI�"�1]�Pҩ�dC��jJ;OH�T�ͪ��4�A�q�%7q�RG�����RT`�tÌ�g�?t�9�T�L���A 3���^3�C�L���K<�\<��i���|�ձ�g}���ݒ�u���|�{���E׽���(�6_������~i��o���UL�`�kod���'�����O�ٽ�N?��֫jɓ	�_��#��%�.[���i�ڵ��Av�<\SUo������ʞ���-ފd���"�"��Y^��������3�՚w��`�Ω�BƁ�*�#��
��U��G��1��3��،�VE\l�#
 �	MLW��Ob�iv����o��p��W��ę��y��Q����[\��B_�p��a�*��S��Ѫ����܋��J�+F!wg�r]���2�Av��2h��u���T�zSz+!3�E�ƉF�Mv�"��S�k����l��\pq�A��A�y|�����&��^[�2x/�_y�̽����p�H�|w�D�y٥~��Ti�l~JX!�+�b��3|f��B�Ѓځ�J��X(�}�|�^S4ܾ��oS���`�9�w�]p�}��B	B����ԅ��},f�h�N7��MG�T���8�����*�1�A��C�:�B��L
��>� ��z��!�PgNF�z�5�/��BH!yJp�r � �o:�}��0rƢB�ا���� �Ck���L���D��i�'jԝ��S#�}�����@[����0T4\��!�PH.FcC� &f���l�#.al<�x�Szbk�q���7џ-��I��k�_����pת���A���U���ҴJ�`b���-f`ưp@YlA�L�L���ߦ��A���М��F��0;
OU��鏸*l�iW+�*!��e��U>j�}�JS_}ۆ��D�74�`���\V���Ev�r*���b�fħ/B����7^jwK��(�����A����l��]�lD��!��wjjD~��,��~6��p���"���x��1o���;{�� �V�X�2@�|1d$��Fܦ��W�T��n��~���$9��kqF��F�Jp��tLY�Q�PȐ	���`�sbyL
�fg������:6�Aq�>2.;����C��f����>\��L��`^��43�Og���"af��:V^HEp���M�.�}̟)��������>W�!��� ����,7���@y%�D���Pqj��+}�@k.�\��[8*B�=g��#��#5*�.�Vm1Ӫ^���F�)m�������J�o�v� 	˷m���"A��?6�a3��J����5fbY ���l�}h��<�yJ�$�˨rf���T!�u��#bɊV���<�3�-y�Gl0�(���ǲXf�����5�V<��K'���ŹP�R���D��`7�����:?T|<�W�/Q{��N/l�i'��s�v��'Qp�P&�fV!.�00u	ȓ�]�*Ԯ+mk����QM�+<�!\�$nϩ�l�"{����V���ee�*��Ci':dS�nx��ց��w��25��:%QG�"�]� ��a!iI�ͷ\{���Z^���q����L!��\S�9�A�]�\�t;�7�<�X�"��^�Ԥ��J�{^��W����j�$�e8]c����0����Q
��$�T���3����9�,�h�Uo�B�/W:�<,p-��@r5�Aq�>~UD��s�y0������rȍ��D��'�(K�����PN`,�\p�)>ܥ��S���H�9���Ws%f���ϸQFh�Z�J��G��1�t$�t.þv%��/�n�S֖c�]x���A�Ơ�w3-�O|zQ0wg��#q�ug�:)��ޚm���Tc8c.�-�<�t���4ɥ��~5��.��F���B-J)�엎����A�b����,�m�wn��nz���(���.A�i�v�O�YCoE�r[��#K{�=�&��S���X^3��L�09����n)�BX���V���t���'�z�hI��}�>��a�ZΣBȠ�#�Z8��~2�p EC�l�7Ox<�]�mm��;��JB�L~g�0f��ҳ�)���w��L�Ψ��<���G�ß����MR�Pz��Em�y
�+!����{)3r�7��e2;
�$k���T?F���K��!�ylQ)�PoE�eU%_@�62�|��oL,Kw=�;��'�dB��G*��ǀ�#���xU���.��2���ot�MBB��m.���|�����xR��؁_�(0ڧ�h��])�=�Ӓ�|�!Q>�nK����A���Uqײ��o�Z�=��៕���Pᩇ��<J&�:*��(ɏޞP��T9;����kJ���)@�ҏ�i�pA}���:.�uR�@�~�Y�,�\�Ȭ���;Q�v�L��N��tMB�6��ej�j�w�cf�f�
�F��g2����X\z�����^	�{^(�Z�؀��\�������&�K	X�D �&�E����5˸ ߟ���+)r���z�����xk���/)�M ^�J:�%�o�5�3���{�ziʸԈ�D��0wB���[ɼ���o�c�{�k�`��b"x�S10Qߞy3�T�x;��)��r5/<��Jc�D�Չ��y�
"0�yu��-J���x�BP��^"�S���c�%��+��3�8��4�������i2��{�S���cέӽ��F�Ң0�ޓ%�j��Z�ߤ_���H����n9� �ײ?���EmÁz:^1�ec�`�>w�nIe�\J5: r�ț\��^�)�6���lMF�{�c�H`E;`�!�?����o�.�w_t@P�� d��q@����`v��oPf�|0:�'k
?��9L ��W�����Ա�`����>/s�������=�4yO`�+f=I�OЌ_�)Oj9�;�ǀ��z�.�L,���L�)�����������K`~�+#cP�������rGO?pe'��������Ƈ�_n���� �(�os�=�����~��_��O8{f2��yd��JC��e{�>w�	&�e�y���hJ����*�4RxH<�W��V�D�eQUI���A�=�@<��.������Z�c���:�8�A��Y�J��,�Z��#S��������L��u9Ԩ�O�����h�̯�W�jF���p�;&p��Z�>J����&:��`cε۬��YR*R���y�U�s�� 7�d'q��`���W�r�WṚ�͚���u$�i��A������yĮ�\�9��H�k�n�9#��N&!I�{��E��w�~ ��+�e��i��O�N-̂P�Ϣ8+�n-�FY�1?�+I�� ���W ��������%5�X�E�<����Kxu�LS!=ɯ��jŐԹzh	��/�O���k-q{�&�no��M%�:�5t7K��:r��[
��2DV��k�ԝ�v�W�ɼ��`}�z�`�<��kf6($�"c&�J��ϗ/c���#�=5���#蕳e���x	��h�a����d�����n`���"��8�z#l���zP��Plcd���u�'kG�!��z��M��H1Q�ڶ�����t�����/�Qcp���np�~c�Ж>�{���I�հljOQ����JyS)kd PM
�UN\y/�kZ����4'h�]��a�B�0f�N"D&]�q�R�U�r�m CZ5Je�[�8�^�.�H�{�?.۬n�����Y����%I���d]���$2��ʛ;Z�����ͣX�y�-sq��i����V
-\F���B����X)gbF�k�t�_�9�s�/{��	��m��E��2\?�o�|��چ�|��e�E{l*�l�b��4��p��~qI��	負���w�oֲz��{��ƑU���O8r�����e�y��T:�d��Og<&���R�J��� ��k� ҹ�9���
�ө[Vy�(������qV��Tb�NR�����U�7@=^X���q񗧳 ���E�A�S�ʑ�fa��x���v�v��Ś!qy��4��,����2OѼ����G��l�Sb�B�w������j��Oq%���̩�턇�!�`56Ώ#C��^j�i���y���'<
��/�zS�>���ᩕ�s�v?�5N�M$0k��"��� ��1ϨP�Ui�V��7l�1<�J�=؊,�b�[�ө��ûR�.W��u��s���qN2�=gs(�z�|��jP��A)kL*�.eA�{�j����K{bW�eזFЧ��rG�h�)�yv�/��ث7��E<�]A�1(���zl��
�:������e��ߥ�qŝݷ�ӧ�O���kE�Ǩ�������3��	!ې�q��om�����_9-��ynL�(��:m�?I��߯G6)�w��<w�CXR�ӈ���WI���]/ 6���Dli��5
:X���f�B����K�����oy���G���x�㙑i�m3|����]~g���O2sWH?Q8����o�b7 w�M�t�G᢮��
�tCd�WJA�)	��#FY�{HP��a��@�>���O������h�R�f��9������<:���Vc��(pZ��;ZN�$��~�����X���a+#�:˟nV"#����q�{��<뼺W�;l��&����5^��JI��NpF�x�3]9�?f�����q~�Em}�C�ɲM�������Z0����o��B���W�04�%�~%|��"�x�r���? �M�$���NZ;\���Y��Op�ٮ#��� S�>8R��Jtoe�gP0� ih�)9/���vƏzxD�F�Ī%0�U�-Mq� P(כ��4I�:A�)���&��n�y8]�P�f�[iY��P)g�b�����I���qm w����,)�Qí���ҿ��w��nq͚����!��s��|%U*����Q��A�=�������W��/U#R+��a��G$ ߲*u��R��Մ+�}+�`���C��PP�92߿6��ۋ�R�	�>�����'�{�p� V[�8V��$f?y�W��Ȏ�wxhɖ{�V,~���NZ�،t��x��fD����)���^�>el����9��Â4b`����۶�z�GU��z�U����;[��G�uOS�!d2�.�o&P�io����������,X�\�e<͆��%�����X��j�����x�?�T5�-pd��`���'���i�n0�΂����Xk�(H�^��ή����8=?��6~�����W���g������:��vq�(��G{�\�5�[l�b����l����R������Q�K�����{�͜���zUrsq�a<�B�w�K�EϢ��4����Iگ}��@�sf<m�@Mqg�,U.;t[tU�nm�P�-p2�v�5$�l�1 ?��Mү+���k뭮�ՙՠ����c�.C9��]Y�0/�Ӕ�]4𒄔���=�����/4Q�����BAe\��fI����I�W�Z�˳>oP��n����6�2�y:I07t}�:0gQf�����b������---���ćNn�H�~���E�g���h����6[���l6aC�����9� ��L�(�t�.
4oJ�-��@���O�+�a��zu��]���zD⅞�0@���3y��3�����v~	�����I�p Xk�sr�VTӿGp�B8���wzJP#���{`�^-��<��|y�	C�u_<1��[��'ةk?.G�_�O%�e�')n�����$?�FJY9U�>?UKJ�i=��A��̻�
��elNk�<� ��w�i�&g|<�����
N*U�y�{�P�>C�LZ�ý$8�k�7rs�e�e���@�/�X6�b�����<;P����� �!��S����$��*K�q��S<PW>[;�A�%|iY����C�Y��Բ�J��y��>d��&��{>���x$Ft�� �=�~��c� Xc�d�=O��%�n�/*��%�S:���p�j5a�m�gr�Wt��Տ�R%�8T%��^�*��π�����|� �Yͣ�\9�NR��/��Xp^�&I˦��oC��s��|��*�B��J��ِ�q
�|R'�W���j�X� F�������F��D~4���xOj�8�n�uxM~dmY�**e܇J�ҍ�*5���jWW�CK
{�|ݥf�5a��j/��͖�YW��n���P9�6�0�/6&�1���h���K�o��F�6I3�N0V�y��ٶ1����	i�}�����t�"թ�H'�b�vKnb��t
��a߅$���;�0�6X�O9�Fͼ}3JD��|5��o���H%DI��Jmk��Z�j���&*�vV>����C�	���d�$��]o�m�'�D>�����OM==�.!N�/$�(a~e��~^[�25n�{05�.4��O�3�
f� �~�=dW���"�?��꿢�w<Ol��!u���.=jk��`�	���n�T����-��Pg6�"A˕+o��^I�&��EH�2�2d��7��!^�[3:����d�J?�c��60���2�&����_sH�,�o$�Q�f9e��L���a�X{y*��3��t3j��G��g��c8��?*ݓ�)&��d�m�\~%���΁C#N��G�0A� �������a� �V�u�wC[n ��.�@��d�!o#�fs�EZ�������#��Eg�}�'A�"��\T��,l\u&�t��aMp�M~�{Da�~2K�2q��'G:@W��r���8�v��N�uDA��q��i0w�TF̱�^T^>�{�����M�¹��cQ5������k��s4g���O���'�WeF��]�[��2K�:a�SI1�&� ʍ�>����r~�R��p���u���qO�FQn�))��b{@\�sjᤶ�j����r�9$f:�u�hB��>�ؠ�VA����5��(Dj�[�^6���-@"���$θǀ���?SyA�M�Ȣ^r�U��O�Q�5oc��"��d/�Ϸ�CE�}���dX3-A2�ҦXv\�x��6�T`��5�6al��x{�leT��0�QpZ]�W�Z�\�����O��e��C`�R[&˂{ٴ��5�Z�?�D ���ð�Z]�	���Te�Q����ɨ9����jM�X��i5FZ��m�1bBƟ�������:�'v�?��?=?�N��f�S3��44���4����I���r��(��Ii ��(H~1��&%fH)[oG�F�V!��D��@�M؛�/���[w`��Mx��<+��ʣ�v�W�t�#f$"n�},���|edA�b��E�>*�⁶gC�Gle�RI��0��C�~�iةw2��D ��W2R�xMF�$4n{���w�����wr�18�.(�e���p��]A:I�%*{@FbF^�EX�n�)��=��@��x �jcPb}Վ0/v�۽������u�H{�71]��/:�Zw-�&��{uR�U�=�98>�����iB���9ܒ��f6Œ�3�n�w�G5[l�5��./�p�������0M��<x�/	H�S�H8t��L��k�볰eY	j�֭�lJ3�\�,ɀ/ćL���:D~�����\��|��y
��9څ�2Q���i���5�:�:�^|�<j�B����9
Q;ƶ׎i�}�N�G4��E�0膖����e�bv(~;Ġ�� � M+�2ؼŴI��0�4��v��7	��V�����Д���H�b��+O��$��J?�|�
.�����]�TWo-ʎ±R8���d7>-���<�����ڮ^ 2�´l�`�\lܡR���T.0�.~��\���Kr�E�J]�G7+��j#�`S�$U�*t�s^Z�a�h�u����Ƕ�d��p蠭7ْ��񭨡��j[|O)8���C����݈��7��u���ژ�]F��@V7бjԳ�A^�8��B��+�F�ߩXN��"�A~@�A�'�ı 9�ei̤��GQ��S�f�F��5���q�ݑv�FVD�q��k�Iҧ &��Ų�U���8��L�'��믩�E���#��c�+��tN��,��OF���7 T9���g
U���=	 ��+�ӝ� ]{]Q�����^��c+E���eJG�Z0�L���D_��Z���2PM���ڿkU���I|���9IK�%/�mBL�1�x��(�m#����h�.��L&��OY���d�_z��p6˱�y���;:�A�+>����q�_Rkf�s=4�3u�b��VE�#)|1���˦5xƯ�݈�g���IJ�i,JO�+���u\��_X��W�#�����JΓ�������!!c�G�]77D[��,(���`
#Z����7�R�G~�%�Ɓ/��ew��6e��c	!]ؒ�%��W�C�X�n�J�:|Ip��~3����z>�����d"Pf�<3)��~-�m<����>q���a�.��0ܘFQҷ�*'F�88Py��hz0~��}1��ftEM �8�9}���|�	��4�N'U8���M|�G(��H:�� ,v�h~�c84?1�k��F�.�s|&?9� ��"�]����no�q��U8 Ff��h���+ bbT�Xe�%�a���G"��x�����FT�py�33fۼ+��'���3�^���+�+��<w����s�����yh����U��\���|ʁ%������'I��>���qvW��ǩ��������v}[\4�6���(�c��\fX�X�O����b����a��F�4�ѕ�9ɿ�~_���S������^��H���(#��㋡���WOH�<�#��&�	Z!�RM��B�S# He���M�l�W�-�����EX�fsr��$t���+5.g�t�.�����F����E��w���?�9B�.D�~O'N�	r���:��+~���i{v-�ѐ�,�-��W�"H�~���_��(	6E5/����V���h{Z����7�2?���h�ۈ/��z��@'��2
1W�U�#���mGq���IL��'��F����g�:����Q�#$�7�!!$�O����c�I ��;t��L�h}�(�3{jz�%��q+�ǒ�TQ��({0C:$���5�Z:z0�y������Zh��k��y��x7�>Z�%P>.8_x��94V��u�+<qF��(��.Qm��t��B%U�&UcI�ۖoF���*�F#�}nӪ -�{�S��CN�����ЎPC���{�o1���>�����o�	͜�$�]�Y����T��+�\����0<��VNs�������O�h��Z{�"��ƃ.��=��:n�;�3�v��z��lf Ğ\�j����S����9������2����ޙ�K�i�j���:
(��}U����w�>=
3��@�a9���}~���{�U(OH��J�n5��(jUMC���L�h���s.L����lrvl�[	Lf��ra��;&ݩʨ�[-;�$�ʚ�P�4�r0я�mC>R��~D�_r�~T.���vS�N�d���Q�&��M��I��9���6�Lx�ێ��0�%����(e0g��i�ςG�|��r��g� ��
P4=�p^����{,�?������'^�*����{
(����*�ۋ�����W,�t�pm��>�����+��⊇��ĺ���f3�'�/j?%M��B}\=��c dU�`H-G|��3���}9�e,lw����M:~�vҋ����x�BBw���3g���^,�?���������[��EF��aP.����);Re�(�ZI)�e�z>^�
#���t��:��rPmt�+��č�+u���E�)�siKJ����aC�l�Q+{��w�)#{^�j�lI�a�X����x�t�s/!���1M!Υy�NE|]<]�`��H��6��L~�I}L4�GG�iF]��w�
���,�f��x��[8�[�DG����Y���Yd����4��%��'��ş�,[�!?��c��v���7����)q4��Ba��׍�8��1$o,:���ď�ܞI�)�\��7�W�k��*F�{���u�|6��Vfm4D���&��@';ɉd.b�@r��J�(7Z�#l�K�'W~Ƞ����^QY�1Ц�r��<mq��-s�+ft����Y����#^/��j9��/��-[�`g���ytl���P��u��}׸��1��,z�m<Zۡ����_�ك¢�Ӂ�i���fbɐ] I肾cS�2�Ƽ���"��cfV���kQW��Y�\4-:3^���]��{\�C���˲6��C�?n_��g���^s�NԮ�(*�0ٞ�$u�H,Ȏ��h�
��jE�I��3i��9`�7#�{����E��l ��+��'�@2y\0we�i��/��F�Տ:>wvT%��{��A�������b��u�J(pY5$��̍a�6�Jn��	r�)���J~�#wZ:M}�����f��RM�|{`��������&9���tV��n�n����M�D����4��"��dpe���K��=c���|�����H�;DT$������l��U�39���:�x.?���}����k��}
)߿~�V�3!�G�Ҿ�����\�c}�W��Z�؏�c��3$����ؑ&`p͇��+/g�kyg��iO�%&�Kzc�������N��5[EI`��On�B,�`�p��dH����:aã���H�]�9��ދg��a������h�co.�14	1��}M�9�u		��z'ǽRlyo*���ރ!����0�2�(6%ORH#u+�,�Zwy�m=_9��pf��Ò�G�.U�٘i6y�V�aT�h��U-B�M�¼�q�Y���<���K�6�:Y��rZ|�.���H�O��Ez�ܵ��f��jV6[� �B{���痸��"�2��Cӧ>1��;)��:�۽��8�!�.��Զ�";��k~�(�],�bkHntw��%�;�{>G\���e �r��Dc����m~Ɂ��GvD�Ds�%X�z�jI�ƫ�3a5��^#�4ܯ�yS3)w�]��qg��o��ob]��>�L��lۏ=�v*!���s�j��K6�RzΘ���p���¾+ 4Cb��:���d̄�����|"���y��ԿYa����y�����m���.�u��1�f'xȜ���8d㽇D�s�z���yR!zю��l7ڔ����Ɯ`�6�cbU@�3yW�<lw�=7_t�S� /�R.bҳ�Dfp�����x�9um�'�7A�I�m��K�r��Ɵ���k[�۹���/�����o�����9�3$����V����:<�7n����8m
�ll�KE5z�aS��R~vK��<��z�]C�LA<ê�'LĦ�Q��r?�Os�����v��V�|�X�6�`x����o�t�ߎ�;���A'�-�~�����Wo�[�9�Ә�;��_6��8w��>B��:��nI�>�q�
ǯE?���.Wzwq�]a��Y���4��k���`/^� ,�J�ݷ�Õs�;	���j�Ѽ�W`����O,˄�����r���.������5[��}��QP�nd%��J������������Z��
��;u{������ӵ*w)Q@x�>��eu�z��-���!�<L
��a+��p�����kx�7���*I�H��P	3d-�8��T|�Q����ݯi�t��b�*^��WP��o�"����QZ3JД,�g�կ`�↉Ok���I�P�K-EA��Ɨ�v��i�jA�|�of��h� ��#��	ZI̚��I c϶k�	���z�9�ܚL�.��.��s�F�qoF>�/�wB��N�}�V�;\�RŤ��0���� =���54x���Ksl�|���lyq�}єb=�ை�� � ,A�==E���9���$b7�/� �vP�1�_q��H����&`��qn�Kz�"Kv�P�>�Մ�`���Q�8�6���S����;�qk\8�7j�$���������x?�4�mIwlIl��>���0t�p&cGJѥ��κ�;.m�MbI���g*%�:�% �՘n܌S䂩Q���Dj���R��|�s�F���ܪ��֯_�pU	%2���&,�ɂ�<�=��j��Px�ok�)>�*a8i���[i?F�xMiB̘tA��=Uk��L��!�{Z��j֥��`d�z�ˀ��Kk�b��W.1dio���B.���F���	șm�eE[� ��Vo�[�:'�ϟzs�D�v4����<��5Ubo�p�ǝl$	b�6���.9+7L��_Y�.��کcL}��s}3�]3��}��e�M�LW	�1I(I�+(31$�?KTG��G�b ���}Ry@|��0E�o=��D����נ��r|�w_s[>/m�p�h|�Y�7FV�l,��� ���`��T�M$(d`���Z��R%c�$]"o��im�������6��bz#h�������{4��~��r��WTGx�0l��j�ym�Q\��[�'{�m���>�׸��P<�un{i��Y%��n X��J�G����|���*e)�����?�Ȍ5V�Nݜ�?s��&�\"<qݍ���۶C�d����qO��!Y���h ]`�"%V�tmXv=���ʠ¹��kE�\>��0}2�8���T@�f�������~"&�(����.B�;e�֌�Z�2���o�\AK'�m�C��)eq��e7"���i�����"�K�����#�"���9� 8���T}�-d�m*���A��3[j"2��K=�p�/�y��B���C[���,ګ1��(E�����a[���&/�����tH��@U</���VA$)��H}���N�Q�����-�e�ڔ_@t^m�O�������Үƞ(F���g�!ԛn�p��YnO�L^�.2Z��`}V��4?aN�$�O{�H�O`�\ݘ�Z��"���N�F \`�z$�جJ3D���J�MK�NEݖ	w��o�Ō�Y;G�u�N���`�s�m(t׀�ɇ���;\���v�r��1�[����A���U�GC�'����0�߹Ix%��E���D�U��Yz܇c�d�	hm1�F'�=
K�三�����.�"􀫿�W��7ږ�@���W���:f^o�~b8�	v�@�x1j��#=�)�q���� ���S�)>��XSϮᄴ��H뜟[Q�$]P����}����֨�4?7y�/��Skh�Nq�#���-�V�ʓyz-g�FHL�$�@:��3�Ǉݖ@�|鱒�pG���Tk5 ��E�B�C�}G[��8��X��O�%�f~Xm�ig��P4Z��8�q�sׂ�xir�kpk,?	�j������UQ�F�"�����al�p�g��^�mf���Nj�Q�oYk˾:`��
*��w�����Z�����C���{���MN}g|qF���<ٔh��� ����HFSr8n�0��'?d@i����	ոH�R���m+U3UK8��0+Vcf���N���0����	ɧ��� �Йԁ�BC��[��f4��6t�����պ[��CYvlP�(_��T�)�T��R�¿�T�9r�)]�j����;v�?Y����轶�Θ�K�ISy;��}J�*ǖ�TECN�>�����T��c���aa9Tv#��pD�e\Ʃ�1��K�Q�1S;��#
��`̱d&S�x��>�4��D����v��|��C����K������C}��D���;����w2���bu�6��}�d�{E��z�sp��LX
������D��t��{S�2�, �-5KW�O-u�(�F�x�<��?z��8T��	:0��<q�.�ha�.������Ő������R)�$�6�e��h������$�RDgJ�[E9|t�a���:N�{���S{�Fo�dѨ�����j�toK��YP%�{�On!*+f���TE&X/�W���L��ڎ~�|Ԫ�jY��<#t>�)Uu�2����j�����3t	 A��9�!�`�s�4b��.�F����w+��U�2A�@�_��A���wZ���\�x�b�G���7��Coߒ~�k��tʁ�&k<Sz��Ιt�bHW��7�aIf�z�k}_,s��Ht\�I������ى̚��/����?V��G��м��O��2IM9��ctN��y[F�|��~+JY7��U�0��-��Qy�ܒ6�L���x���q�:K�j�!p�4�߫Ѡ�Ü�zu�s��0[������p�QJh���ȳӇ�\��)�t��X�����B���b�t�2�ֶ��)�rd�}����Q;jk38�a�`��y!K��{�ۨ(��ж�=Y���x`o�+�!V�Fi�ΈO�*�kw2h�i��~�}���S���y���"��K7xs����$[0o�\�Ȏ�Z�x䬀�,״��I�=�sD��B4�(�`6��&�?{��n�)�<�%/%�� �GB��\�:Ę�����M��`!s�K�m�(N���+!�+�G)�k�_�Se?P7�_�+����X���i[�����~"(|�]��0��n4���*i1��H��S���]�.�����u�u����#wF��\�b��_ �����6S@���Z ��`�6k��,c�?�����X͟`�x��mG��w��X� t�`69��j��ԹF�탒 �К-��P}�n5��mT�2��ñ�;��^�������~�ar��h<!G�>-��J�u&�wJ>G����F�}8����%|�r��bTM��ts{� ���_�����Y��9)B�7 ~,ٱ�Q\�xT���!
ک�@���{���O��2�(.l5dH�IQU�
��|����u��[.��<�@��'�`7D�J�+�C�{�m�H���J3O�ñB\���%j���Y�V�3V[{Q��I���(��F��A^�\��?�7��n����H�{]p��Q����������f�,�ܦ�Dh��7�`�%.7���vOP�V奶j+Jf�;e)���G�)Te�}-���"��YP�j}��L�$*�f9��'Q(+N߳�W��p�g^����9��4�?���o�/��JAKE|���"O�� Et�yL�#�|<m��@k�v�v?���pf[xL24
�`{9����,��  '�����3rN4(�����	����5��.Z!���/��S���fC�u�#T0͙&��D�j�d�18�.�>og�(�#���TL٦\DD��
7�r���2�9H�_�^7��y�gV�%�`�����ޒ���T���EdI`�l\�|x�_�����W��!l8�O ��fԷX�u��������n���h��-\��q�4\� ��
2Q;�sۊ���l�,��ڕ�q�)�cp��T%�FqA��7��_K���(�P���\ �u(8G�ox��'�AJ�%E�2z�i�[3ԿӒ� +���[faG�%��w��W�v*jcYA��/'��p��&��L�x�F
ێ�մ��~����bX�:T�H.����R�0���CӼ�g�Dp���EO)��`��w@�#:�:��]z]j������Pq��Y��Nvѯ� M�N�9�J���0i(��Qrz�����k�%��q9��� 題�T7u�kE��C���/،)��=b�|�K "a��z��N���vtJ�c��;��˝pS�g��n�z��?�L,G�G�e�m�/7�	�D�ky��''�a4<�p��U+�vLB�?(�kk�����9��r�������lyeV�S���WB6������@y�#�}̼��P w����y�r��1���>$[D0���j�%���Iegp����nY���;����!)��P��@N���eU��h�);IV+�׳�� x8
2 
����T�/m`I�Qp<�;��	�+����ͮ�gR�l�#�1o�[rto��ʋʯ(��1��;���֑��;|�!����_�[�3��W3�P� %����V�G�
���ҠNg�gļ{�Ij�Nl�@�R�@�'!<�ye۠�R�r�5���
���4-.q:�E�����V7bI��{2z��$CҘ�/z�u�-Fcw��;�#c:��0Úǩ��t�����dCb��;�����"��.h9moKǳIЯ��93�����K����.���r�r&�[	7~g�#.�8j9��9d@��8z�2E�8�tf��wN�,x$d�X�l�۷na]�rK�Q[�~k��o�g�䕓�~��:v ����r;x�佘Y�$
�B�|�勉!�d�����ha�J��DLvT.��ctɉ� 	�Ƨ��.���V0j�	@���"�'�A:q��z�{�lO)��§l�W3��?v�5?�qg�s�B6�ɰ������x?{wͰ[�r����ʬvǭGu�O��5�DvE�)8���voo��B?q2�g񤅭�k��%)�V�v�vq�:�����-���|��M�E֞��&P��[�&-�n�GN����-½�'k�&�a
ǚV��W����mC�r�eW�{�W��%(�zϺ�_)��qE�� �k�8R���C�A���ث*/��ܘ�Z1�+sA���.g!:L/�1+E�r�ۯ[ްwJ�)N]ՈsI#����
�؏��J��`Vj�H�,.��~�Ⅽ�F~�0�1�@�)x��	_{���Z<g���������
�ξ��A3v�t�3>$^�oJ�u.��ڏ � ק�]��/M~zV��b�Q��P�G[��Pve�|A~'��sy���5h6�&|tXUꖘc*	�W;�ˎ�O�O)���<�����W�4��;!�����F��9��rě�y��z���W�k;Nb�u9�-7�B����+��Jt����,'��uЭ���nL.�O���$�-�Ad��])&��� ޷.��:נ�i�����@����Rj���DS�./�Ҕ���I���`U,F�ĳ�;�ER_��םt����q�:��-�l�4/m��� X��8}�!�!�p{�_P���F4u�m(�BR�ﺐ_��������6��[ר�Ҽ�C����n)���j��4P�!k�?�)Z����c������+����3�;R2�Q�"��{mT6?�At�2~)��@|˞;W��oL�!�[u�7ȸX�j�c�S��pj�����	Yo;/M�qǉ:�_|���[�F@�ݞ?b4�@��i�5���m��?���!R2��� �6����������ʣ>��X�F�Ѷ���!�zl��\Ț�'fa�)�f�Q�+I�v���s5ޛ�wZԛZ3_�N�(J����n�zƶ=���B�h(�w���c�w�
�Sw���j�c�Ρ�G]�ֺ$�fʫ�;Q_?�v�G
�Demr���{����N�����Jݪ�Y��F�Dڷ�W����V���%��e,�Z�ڭ�jB��#����@Q��Hp��ʮ����	-�c瑔�	��9�)��1\���PW�On�\�*���X��J
���7��]Զ������b����W^�9rS������:�w�{��e�T����0��X(H]��6�GJ<�}�V�g��P�?ˊ�<��A{n$��� B��|єlu�og��[�+W��]�C��U���M⌑v?�%���t��Z���7e�v�=�5�+�Jʩ�7�$���S�.%�12a��$���Պ��O)1�4�h���TH�k[CD n�<ָ*�D��ϩd���ѬF��/5��nS�F-��J`o�kd�x?����G��͕�����(�$�!�18�:��3�^��YHiq�'����d��o'�=#����V允��q�|��Po�
gH	���G��]���L�>&���q�����҉5�\^�����%�Fڽ�~�RǬz��aܺ!�ĢS�a�����|�L��QB�:�"fH��f�2�͍�k�@��{�g���������H�1���
�����lͩĿs~���|�<����"Y������Kщ�:�0ٍ��ٜi�`�s����+v������7�	������,��>�eg��y>��q��r0�'M��c�i-��7��tbβ?�-�rj	��V��ɡ?���z��Dg?Q�
�tz�c�[B3�8<ϴ�4�=i1��nUe	�_�T�6y�gn������r�a�;��;��Q�m ��D���h��O����3��<!��7M�W݊d�E�(>J����.�F�;�CDNd}���0���V�_�ٸp�'f�Za4����Y�������(��݌�������c���+Qq	��gbl kM����8x��9Gg3��V�X�ɭd�~��6x�)���[���9�U<m汏M���85�X.�.K��f�5�X�:	��E�U�6�����iұ�Ԑa�YS�\�`�&˭33Q�fkd����̩�:�:A��\��l�I�vOAjk(R+|���d�V�d;LSQx�`��Mȃw���5���ۭ+���2�Xj��F�xa����lo+�s�����#�X6��f�o��ka���R�z(�h�Z��Gt��٥�&3�#r5�\IV�/\��e�ݼ+ITR��+�k1�k��8,��x�/�W�;��M��f��>0y��{��q���oMG��l �,�X�*�;������'�뚄r�+�>�X�qS�k���5ؗir�v)M�E@F<w�o�,��X���+uk✅�bm2�d���~��ڏ���V9@�p�}�g���MR�N.�i�}�h���'n�'r�Н�W�9U�F�ul�j�����c;Q��� c^7!��׸�.
���5tɝ��
) 1�V`F�Ռ�ϼ
6鉌��ls|'Q~���'��h�ޜO^mr�<F��<.�P2�_��;W�nݰ�!{S�p�u���L����ҟ�(1���4��Xo&�Xr�`���2�6m�X�Wk��=�&�4Z&T�h`.�ڪ� #��_���Ӕ?^��/wf�O8^P�8�p�ɚ�(qĔ�����+� �"��W��g���A��վ�^ ��#{�i�s�$�g�'k ޵K��Q>-D��^Ϥ��9���Hp���zz(ދq���k��h_[���YQbi���"V�X�@ݠ�B�w��.r5����Ю׿խ��!���\Q�ihyW,�i�oŧ����G��f�,/��+O�}O+pW#�CƧy��9;@�М�X�=��MO~�������X���	�'SZm2Q�35��]����Hiv�??���VO�� r�.���`O��4�5�]����0F}#����y����W2v3U
��(0���sfV�g��aY�-�g?;��9��J�L�ͱD�"���j��$���t����F�T�<�N�2`P����&y��`�Ɉ�j�AR�X��r��pU���Bc<���P�����v�	w^��_A"��7ۃ.R�)z^p�Z���ͧ!н��u�LSm���k3�bѠ�枘l;!����G墚�W�ReӅ��>��L����"6f֏3�N�z������L;�Ȏ�1qV}H�ime��]2�9�5��ދ	�.����Z�8�B9��׉���U��.����W���� �}Ń`-
�%Q��]}�KJ�*./QL?�e}5�/�Q��w[���y=������@��rѳ{�A��ܹ%��_���~_����Φ��g�c�
[e���gGA�����ϴ���.5~�gӝڸ(4��Ԣ'Y�o���Wc��/�ܧ5��r��q�R�^��!;B1s�e���zM����b�hi�=.�g7�+����0�?��`�X��]?�&���%���U�2쥊פ�;��ܽ�oXW_�3�a��ъf���G3�U>/��,j�.H�OHf�y��	%���8V�h|d���u_��}�%���|��O�[�D�#��y&������z_�'�Ɣ���4�Y�H��E�
�U�;�2�j�5Z�����|]�L����6>��Bm��ϡH��>C���anqz{l,�-q�h��R���6�X���'�f�H���bz���	sA��GS�}�)6�X����ޝ��WV�h�/�����?�%��rq�,�dn��/J�e��,SkB fC!���k�;�)�A[NcK���PL�J$]�?�I@����%�8���W��X��(��y�lN�(fs�I�¼�(6|�[doU��*
"���^rQYСHkY+�'�V���
e7M��,�6�b��z�.�e����m���f#����?7�rE���l��Q<?#G���N=g�_�FO�A���v��Fё[���������}�a�C[e�&���wgB�i!6�sK�V����R�ny-sD`)�5���]kZ���HZ���,�}�eO�t��^��s[�4�+$���y��
�W.yC'_���fiI��4W��RA�g�I���J�*�~N�ZE����Sb*2l}��̃&Lt�_ۂij"+�A1�(�@�5�k�Mkp�<���p珻K�B`�v�
��C��t���6n��eJ�>�Z��H9d}�*���^J?��DmU�x_�R�t�xX;��{�z�����F<��\��$�W]fz�\b�D33b�ޞq$�ד�>|��=�1��J����\FR�@��0�T`�:��]U�_�[�KQ��529$	z]��"EĜM�����rx�,ǒ@w��D�(~��'�52������G|$.��1'�6��1��/�|w�6�A�;� ё΁�p�wA;�e�jT����Ԙ'�����ť��m�iH�ϐ2^qQd]��,->m��1ZS��US!�uόTZ���NM���,5���1����5�������){cmQ@z>��5��I��{�ɋ�-d�P K�.�~���#L�>@K6��,�ѻ����^W�����}�~��n72�Ǭ��;ɺdO�\�nn��g�,�@�kиU�.�mA�A��ld����I�t��H��IJ��D]^x�mŬ�vE�^Y#���0�>s�b�!��]8[j�(V#�Nwtҙ]���um̺NW��C���U�u�Y`��r�����[6#������:��z�pq��nh>kGC�ZjF�d�Z=����������p�1iX6`w�O�g�ǣК1!�����<�JR�<����{FG۹L�q��qK�i	ה�E��P���K1u6�Vr���?���ޟ���]?�5xi
EO���ܜ���;��m��LXs��Q�� �(|�{oH���i��Y*d:-����ׁi/0�ZU3�ǭ��+����G��ˇG	6��P&5�S��2w�*avu
4�^�L��4����ij�D;h�J�^x䝃w �u)$���-�f��q`��SOV���\K��t*��N��Ha��*s @��E����z4vF�y�B��/ �\d�g�¨��t�H4��b|4��}���-���t�����3���̔:/bw��ϛ?MH�\��V�3���TR*uY�o�ҧ~IJ�F��g�1	��$��$�Z?k��BR˪F����u������c^\�.�Ac\��FT��b�w��r���LLw����Q�6�҈D�S쳆vP8�T��bim�b�NJdR��2��K���vhxf�P��sq��y?s�jz].6����8h]��;����T��y�l>"�D���S����Be'*ն2S�jj%߽gl�ʅ ���;|��-�z��a�=aA���Pg���(����b2�������C�
z<�rf�F�V�`���d{|��ڱՐ��֟)�7�����J���d�`�hob5��6�l��ٌ�ѺQ�QT����Kk��_G�6ed�D7����x'��[�N��(|�E
�I�$���`�1t�cx�ю�$��{UX5"�Ž2��A�AW�Y�O�ぃ�!�L�K
?)���i+Q�:�F�E��⵰��5v,��T	�8DE���E�q:U�������g,�>�˃`���3�õ���5�F_���3�fn���e�$-W��m���D��܆�T���\Te�=)�	�]@����e.�����w��?����P!t��]�q�V�P�]��9����Hvm6��Y�8X�Q<�>��z��]�k�d����¼OڮMJ&R���ؖ&YU�D�<�������&�����UV���a�Uk\4"Pꤻt羖<��r�|^�j#'���ٍ|l�&JP~���kF-�~i�U�s�Q���]�h����rP��@˂a)Ƅ�D9*�?�e�u� �e�ݵ1r�L�� y,�-uz�+Jpe�:��\���{e/
�^G�?��{f=�Sq�l�ǫ�{���K�G�R�����e�j��#�K�⚛E��"N&�H�-}��A v�&\���:��*T~?�8KS�3�a~Ɲ�H�_\�>��7-��œ��nX7������D�S�GA��W�h�QMf˴X�k�#X��>�����������+UniM����h�R�{n�� ��)�X��I� �@�$��ѩw�Q�ףE$��9�w��L�j)L5�_�y��.�a��ԕ�@)��x{����4�\�
���ғ{ya�����_��l�nU���k@�g+l��c�/-F �f�`�`���'|�h�Ask�oMg��{14_��r=m:ڤ�?����cA�A��g���b����9����;zL��HA*̳�g�(J'㉃P�����!������ �hRmo��~P�25�����ת���W��^�� ������F>�2<}�����gk�RQH�B�	^��_3ȩvhr3��P�c;; ���B��E^��_K��ʉ��lD�<�\.�0�II��i_�H�n�)��|���8�J�Sc�^�T�O����a&<aW��AH�҃���L���?� �SӴc�u���i��YW|�q(r�ٰ^F�/���o�����~�4��د�>Qf��eIV�w���jPU�Ҷ}=�����r"�S��	v�gm���*T�6��C��Ch�Z�w�ó|���D�\c���y�h4��_��\�A�(U1���f�������f�,�S�صΗΎR��s#*F`�����Q+6�{h�Wއ%�c�t�1�O	�Vj�R������~�������P�i�i��V����ve}�B���K�!ͨ�h���Ւ�K�z8�l�M>�N���1�Կ,!����`�,sL��\�f6xo��z�Ƴ[D��hKP3�V�
E9 9`B�RӤa���W\=�8N���)�'юZL��9A�M�,e�ݺq��Espy��*�́R�������v�ձ�C���g�MRm���xQf�~p!��lZ���>���C\N��d�����ް���a�x���X���aԘ��8Le�#��t�	�w�q��S�7+���:��5B����c2r������}��cC��U*�3��Ͼ �3�t�����#�	^���#J\�5ز��K6����,���m��`�pCpS��⇾ͫe5�����Q��^�[�yRs���EJ�I����0������Т�[����wX�IqW�S�;���6�څMw\AD/p�ə?�b]����1v�?�,��q�{sb	/����g��9tǞ�E�u�pl�6��� ���4{���x�D��pdvNG*�1>B���R�%Ǿ�q,݆���5o�k51��uO���.|"�-��B�	���xR��J)-y����f��Iy�- �Ϝ��.�T�!����,>=�i~i��ݼ��Q^����gS��[
GX�H���0��[ �ZI@�.��y�lĒ��ir��n���o�X���Y8�s��`d3����<�|�J�lb�<u��vP.�U~pk��}�T�y�&�A�|Fx�g����4c3�^qM���
�����?��S���ɩ�<�~���U����J��bo�=6�>U !2KP� v�B��6V�W��9�}o�'�q�R���K`g��:N�KB�6�@8{@D�G:^��U�7nS��|W�b�?��5,h/���b�W�w~�y��Fd$x_��L4� �N��1[�� O��w����MΩ)��~8<W�8K�E_߁�D�S��{�1��mv���߽�7J����^,o1+�7�gr�w3.�{=�����5�GE�wx��d6e6�=�خa�:��L��!��	\G�׿�e��XO[/3���!T��&k��?��5d�76�4�Q�jk��L�P v�� TP�o5�Z�s�Q`�-vg0���8m��k!!�y�� 2�M_���r�c���zB��@ܜ����Xd�04����Sԙ�C�n)cP��a�}�c	�R���iR��e�C���6����HA�|)
�8��Q�1�.M�M)�����^��ۻ�,�= ��xU���h��W��u�:,��,��[�0 Ȑp���A�F�o>�Wo{�Q�����4����v[���6Fґa�A�-�R�E���Iw���2Kj�INN�rN�X�Au�>�6<�S���V�7_ܥ�k�<ݝ�~�<�Ts��8�)O{��G|�yn��@߰a�4ǘ�Y}�$Aq��{�����>�=���=@S�8�&&>��#�zPPJ��am������=��c��߹��4�+ᛠÌ���<��m�"������ĳ듘��{�
"7(Yw�%�^2���.7��H�4��^�P��`2'�����˯Qq�fA,ħ��E3GU�_@��=�ز��C�h���U8�9}�ޮ�p�R� e'+S)��kE^�Q��s�	�z�+΢�QF��>�V�jX� u%��DW<uŷ�7~��툋�T"Uv�8�C�P4l`@�mn^a� d�������w?1�� 971��'�T�<s�z��9��6Sc	��B5_�p^��λ�1BO��]9�)�+�%ȵŸ̜/j��W�S����W�qZT:\2��'v�}�9�x^�*���6�P�mLI��柵��%�se�C��^n���+���H��wo���|��7B#2yr�DSY�h�p��v����e���/�zh���-���^Q��]��T�:��y=IN��,l���N��"PT{����&Ï��gTq�]ώ�&���i��3Lt��
�ԂD//�tl�½[�r�s���Sv0
���O��Z!�X= ʘ����S��Xd*��q9�(�L3�{t=AMc,�a��$˴lS����>ENr�|�F�Bo���[�G %@!�s/��:�	�j�	HU�|������!}�:8�S���N7���.�c����8Ģ�纊e	���I1�D0���7�$6.���(@J�߅�ͳj�y�D�;�	É��rq���-U�7^��)�N�墕.儴c�xbzV:���P$9��U����4O~%O�6I�'��}�&�
�9���R&��we�r糈���N���%����n��(��M�m�ߙ�������+��w�g����AI��	]R�����O�
d��p��Fr�����'$�C�W:|�b�\r�剁�X�y��<q�z�20�NB�
0cs���� �U�Q�%�n���[ID~{4��~M���1L��|C)�IQ���xϮ-K�i�������]f!jq��3�(ݴ�� �+�C��:���`�x�4Ӱ�� 5z_�L/��*.c��D8�E���us���{�dcw]ZV����	����k��kn��GJw���VH��5�)
����Ӳ�6��P�/��25V�(fξf�{F> ��#�������;ރ�����)�h�Q;��~� �:ޞ����������i����[S��uW�ރ���h�Z+҃:�Tr/�Ðh�)����E\��T��)bDM$\�����-�qYZ�n䋱��a�'YV� ���.��^����ю�W�*%h�����bh�G��%��O�~tjX��^�Q��0E*-=�63Tߞ���
�$�`��$U��O>�v��7�_:�Tue�����g���k��'s����H�7-����"@��2������� �q2Pq�i rE[��XPo��c>=�p	
�}v�I0�t*Ϫ�Y��ik�e̝Z��f�TQE��^ac"u�j֒�C�䦈�ph��ԬJ_l��؋h�M~�2����ň���ѭ�����J��p������\6�T����2/�ϙ@<!��ޓj:�N�����u[J>q��5,�א~�^�%���~�<V�]�'Z¸:w�2�VS
Ү+�����r�1& e��*�Q�$�tb��p������tg!��}���I]:��T�<
��z0�1�/�V�{��4�����(p,9�%��ܨ���S~ L�ҬL]v����%ء$�Lm�f�i�����!%���٤��,'R<��>��Z���I�#���=�ҷ��o}S�4%[��Ǝc'�-��eb��$ѕ]�ZK��H;�LC��GؘT'��߷���2g�����MvZy��t.u�I6�f����IΡH�� �b��	��sЫ�<C�����z�w6t�`s5�]�i���:!�Y�ؾX�C�/6�uC5~C1���2٭�t��AWz�$L���W��tM��Ae�T�QVC��(��N>(������C���Ƕ��A�zC���j�+��f˭\o[.]�c��pr���0g���O#"0��/H�o�#�������Wޘ}��˛Ҧ�����6�zw�cAG�������?���J	C�ri�HjAr�	�N��]���@/� �)�<t��Ϟ�.�v/R��{���;�a\�D���橬FK�e��0�
��XN_R����f9Z�����B�$�pW�T�U�`Q���g:0�潗B�<J<z��U���*Cn�n�xX��q�(j���ڽ�i�y����� �1�k��>b1��7����ƈ8��>��+g��Э���G�� �ۯ�7\�U�[V��W�ُRc��b��u
�<�i��W�v��`Yn��6U���!w��{;ZL�xٚ�Rӛ�spNr�b��������\x9���43Q��X!�&��0L�_� �� 95�(|�5��{���5z8��z�y�8I�𜁆J�E��J1U:��	��n�yg��^��C���{}ss�ˀ�mԟ�[�^�3�S��)�}@�d<8)��`Q���鷞�L���tڽ��|C��E�
4�DP�-4.��Iz:�C��c�j�Zj����QU~� ֜`5y�y��@���� l���:��U���͘��>R[H���Z�4dΔ�Pg1<���=9�p��b9��*�rl��6��'4�����UM���$ ͙a�����ݠv�^
������e�`�Ӝ�� ߄�=�d�p�u��z��j��3�5�4Y��&��r�������?��V�f�\�Ip�(�lO[�䵿ҕ`��P��5��q}Aep��f����T���%'cد#|�p�x_p�!�YA�D�w0�^|*7k����ȳ�<�I��6��3�s{c�J����ͫp��D�G��~�$|�a<䀀R���4*�W%�//���/�S�;������6-���qlz�^۪"fz4-�uy�>�Ԝ4��,��<!rv�1�����p�.�u�;�E�Q����hFγ�"{�0���� f�qN��}� �
������X��k��曆�Y
��(�N��	�m��~W"�7;�:D��C,�Vu ��/:���*�-�M+�X��N�ǉ.�����j���A|#���F;�6��2����lVȶ�����ԶU&3�i��S�4��O}�eV۞ ���׀S# MoP����cmj�%��Ę��OQ�I�ў� ��̣!�3��Zx�ZU��a�$q����MJ2һ��*$�@mԺ�D����#s(��6�3���`��ભ%.�ƶ�A�6sHҬ ���ۨ��ȕ,�N:�)�f'�	���lR�2u�HPk����{����[�+L[��V�T�9��R���Haz_Tq�~��z�b�qq>��t��<:��HPmph� �S���i���4�j[�z����&Aq���3m�?�m8G�B�s�y���0�W1sc�lL�Pxs�(I�n������-��� c=\�(t(a3�ޒ���f��ڊ��0�v��ź�KcW^~�������qϥ,?�j�b�0P�5�պ���������;��:�q��CC"�ׄ�[��!�`�En��Q�-{��
�������G��,��9V�0��~��	L����p�^�2
a#iL�E1�4���Wm���N1q� ���?�,;��4��G�L���alY���Շ�ݬ��!D�i�G=� xt~/Hz�dsY��`F��8я]m��~����u�n���&2ޣ��(��[�[����<�߂��g�/:��;��.�v�߉�%+�v_Y������=�>ˬ�ˀI��ƞ�d���g69E@lq�|��Tt+�qvdЕ>E9\���X�>�8c�U%C��W�� VFZJ��'J;4���m`j� P�S�Ud�����;d�z�����j�j�`42�L�yI����j]�;5A�K)�6>� ۹`�pTBR��4��.y������R�ſ�㸁��`��/�@/y�"n�k�Mb����e#�z/�L�V����-�T�gY�m)���V>T�J�g1��F%�hM��kG`^g��PP���� �q�O�xç��F� ��§��b^��*�!
�{�U�?�%R���{@����L��������(F;�5��p��R0���HV}K����"�w��Ik���v�E�4<4� �Q�mM���B���P���G�ʳ�{��VU������Vy��:G:ܤ�$��� �tkfc�m���ܭ+1�L��W	���@��2�ǤAN�BK���J�In�t@���4EB�z%	[>�'dA���z�q��ǝȂ�f������n�����ƋB?��}X�����-���寘��5gy ��z�P3;��F+uV��[VaT��٬\B|��3�&��%)g�p���S�*�t�u�,s�ZA\N?ڽ:���šw4kx0���1�`2}M ��蕏僺pj�&��Hy��#�X^��_X��!f՛'c^h�R_�W��L��c.{)���2�1��׵��N�^��z�7�+�?:��T�>8�0\�U,�4[��]����x�%�F�^}V$�蛻�L��/�4�c$a�|���6s&��o�ů�:B'~��`P�V[c���̔ �*^���`	8)��7�A�I,���ig����Ԧ�3�mu�c)�o��E\)�Z�� �� � ���;�K����9���m&�ŞjWNƤ�T{����FF�`G��AZ���Dн�<�?x�����taI)��뼉G�*����N�b}� |�I��g���Q�T��	ߥ��Zv�%�w�P�ˠ��Lhd��6��;�7�o� C�m�lc�uy���C7#(h6���4g��@k�/Ǝ��Q�V�S���-~ha=Sw�$�.��>�n�K`��(9vuo�͓��JZXMOnZ��b��,�yh�1��;�*��W�q**P�
�]���@��n��')�؅9v��Z��]8{��R�$4��*�ͦ7~��=�P�D���h��8�k̓اRi�$ظ�ٽ��.���HǼ��1xOO];��V  �M��D!�h.����5:;u<a�SZ&#�<�Ǌ�d<��|�v�>ϗ���|���*��e`b�MɌ��Ϛ���S/�ʡB���n�F�c;[����K���"|K\�nw�-�'m�3�N��yp����#~��?����R���rb��ӈ$�I\z��yq�@dRSv��Q��^�E��S��q�"���>�/��g���� �F;%��m�.#g$j�&��&���d) Df�б�&�Z7�7AL���!`rm�^Wd۱����v���Aq����� ���rwDҿf�{�l��Pnq<���q�t�5IO�z�i4'b���u/�-꼧�[n������ҕ��j��0XH�%�o7���>Aj�C,M��sT�6�~�l�bj�=ŗܩDDg�Z9Q@f_�Q���-���y�����pm�n>-9�E�������䇎����V�!Rzq<s4SI,�*9�V���q-ju�e���C-h�4r��j3�ΰQ6�l��'� ��$�?�����_I�l�U65��xGEw7³��7	�D�kCnuk%���z͑��=�W���2��E�8M��q")�S�e��D[���4��� ��*ӐFcb�y�a>��!�2���%��T9׽3&V#�oD�|�Is��qݲ�C9J�U
��N�6�Y�֏P��0,7#�<��K�J��>L���v�ǯ��Ph~/��O���6{����6�Yy��ϱ4�zr��Pq����K��4���$�^j]��޿*ʺ	�#�����_QҺYv���{�mcϞ,�o)Oy7^x'�>��#Rq���݈4�5$�::Z?l�52���z%���E�j����1�SK�l��r�8��gpV����q�x�-Û�kʓ�����&�}̹���0hz"O�:�֑y�V�z	ɢ�4��M	�4���dB�[�D%|��X�?Dh�\*v��:͎�l.��?�Z=K�=m5�������V��Qo��_��W���Y���s�mn�#~{��ٜ�)�])I������-@w�ǰ�Ez�Vfs�)z�<��)ȭ�L�\{�[��sĒ�E������݁|�H'P"�Tlmʈp �p'L�))��׬y:,�͙j!�� k��y��Xseyp�k`xM�IOo'�ėSJ��3�����2�����:��>Gς��_�]�0����y�?��E�x8�V�0v� 89�v������� D&�B�_�������î>~���7���*SqS(&���R���s�sr]��n_f�}9L�̚y�,�H��h)!Ӹd3�6�N�4t�]J�ĕ��Q���\�zʴLò��6�dԜ�'6��M�Ph����;�7^+��ʕH&�!Z�گ�i>�d¿��5���
���2Hy����Op��x���UY����]�1�H�� r�����h��
���R���w:��b�ʘ��  gc�'w�	W�&xy�n'|��?�67�3_TE����̈́W�y�g=-��27�M|��4V����!�h�mMS�`j�ûR��I�1RA���a���"���1�
����i��WԪGs.���N�n���^����6nhѼ�X����lu`�T�ȫܶM��̗�M=�Utߟ�7������(*Q��s`i�ݱ�}X	�,���{/r��֛� A|��IB�8@���6��z��b$��M�I�3�~C &j\��G�?+��ZT퇯.� �����.��N`[�"���h쮪$�	���{|����k�/�-x\La]6��9�S)�?8Ïh!*H����۟#�fu�M�?rǼF��,0'|Ծ��̎�; ��|b�
-i#n3	'��նMٮ8�7��C�0`Ս�H|ʇ�08�{�c�N	!M%y���`fJA���$���/��Q?�9�Zq/��|����T���┓ ��O�ޞ��x�>7��(s�Q��b�{�c��W�j�T���qv�A�?ژ>5�����G����<���#�f�L�O?�4��bj/�.���u�g�ʂ -aݔ���V)7�b��n�1��d��ð�N�2˟�S}���0q�*-ri��Q�#Wyn'����1T��j�� Wx;f��]�b<�B�!�C��� ~� h��s�H��U��$r�>к�l� �V�h@�%��,�iȗ�������V��i2B� �R�fE�AT���e�V�����QY�)N���7����0`.f>{�R�?�I�4�1Ii�+�KKy'��a����=�B�p7�����d����Fī�2��є-��%��1�+��n'Wx^3�=o8�YK��qƜ�Rݟ��#XgI���o�������:�p�y+��:�;�0�Og
��[�PP���m�|��0���z�SFM���4�;Or�V!�|�l�b�b����>C��MfF�X����s���}*��^fPV��6hh<)�bbf`���f{�n�ܽ��MD�Ga ��`�!@f��ا�:�d�R�vAc9�=G3���3��Fz�����вU�Qj�:�<�{�̷\��Λ	�}����� G�F������ͼ^Y�����w 4dc�sCW�9�mƇ"�$�`U'uZD=��$ņ��Eٷ%l�Jw,���|$%��� }-8掽�����)�#csD�t��e�G`��E�������f���m �+P)��a�ƻ���*�5Gv_v�� �B��k���'G�%!�B��:�>%���q��v�R1�����_K�s���ij�o��y�f��KP"�J��aQ��������	ȃ^�^�|�1���"$�����u8�.[U^��?���]��/��J�ˑS�jRĀJ��ߵO��k�@%��qx�؜
��f�$�"�C�	�sbn{g�}_�3�s*G>f��Oq[p���oӅ��BK���pL;����R|s�^'�sn˯¡ڂl���}A@)�6�aث�)̡���FTuq�Q�T��Gӛ�}ދ��rk4 ?"�=���8�Y#]=�w��0eN�H���^nV$ C҆g��p�9>G��� ��s�6N������M*�VcZ��`T�;em\���ās��I&a�1��:C\�Ī�w7'�8�Ό�����$�^����Z��́�����fO{|�����ѭ�A����	[/���TvJ���:��Ty��������,5�����nր�w���
R?����`^_���EȒA���9r���B�J8=�2O�uvl��ޖa;:���=2_	Q5���|\�#����y�
�O}yY>�Q
'�������ٍ♭�_���7�9���wdc��=7�M_�ۙ_B���$�~ؠݲ�dIjJ�����v)�${��H#SoR��Q�9R)[@=l-T�u������^�}pa�z�1���S~ӌ�eUCHp^��,����o�����ՉLT��4ѐ���<w�&��D�[�o�12b!�[��rE����!:�H�X#t�@�N4j�f=�0s���FLm���/��� �Y�X�fcv��0�2w�jp�h�y����o��3�D���n+�(��Un�������Eq� �����m;Ԏ6�X��ݠ��U�F�%�����D���7V,Am�F�pg-��5�qO����q�}���X�7Y�d$�:��ɹ�ȣf��$	��p�TA��l}�Q�]�'O�dy�vRd��3�s��_�X_"���=:�O�V�b��9�ߕ�_�O�'9����v�R^� �֨�����ĺ���	8�M��_dݟy�*m'�Õ����M.������'
�s�fu���%�h�hwz�Y��s�l����x��>f��8YG$�vߠ�*o��8د�����U��*�cr��[l NʨͣB��*�Gh�΀��
2O	��E5�6�l�
�`(dt5["�E�!�\���]�c���F�cP�����0j/��*+*��'n��wF�<D�1y� ��V7�JAIsެ>�3�c�X�!O���/�9���l��5���w�֯��tŗR�r��[���
�z>�'��}lRA���-9b&��KO���V\��O$ǃ�!�a���V0�#�:X?�f�o�$Vd�}LO_�
�UцMה���j�A^�3ii�V���n�;����z���ߏ����2E�N���׌)�ya��'!��H��7 8���tg���Z��F%D(�Lꩺ���P��s����Z����W�U�����C�fm�j�V�͟E���6}�sk��x�u��V�sX��Dc�����o
uX�!����'���qq]l��E.8��V��@�V^�B��:$�#6=������J�o���>��!P�IT)�'���zɬ˝샧�6��0�+�,����>�Ta�ؼAO%�Hn/b��U�#�!h�L08�2�j_��f�A���Tc曋�Zв�ڔ|��k�
P����VQw���?��<Phq�[�5�9�;]Ը�)�Ѐ�|Y) �M�b�_AyX��&&�tF��}.T�7�7�/kG��V�n���3tv���7����𴬖�s�L�<�����ZR�*��o9֊fg_RsO��d����ܸ%���-�*n�yN�l���f��8e����E7b=?J�4��9�N@�as�������	s$�N٧�l��1n?����L��\.�~tc��M׾�����	.eJ&nCW��s�^��*{�N�ӈ��d��"N���ѹoQ#e���m����2�q�����c�\�w��&t��ɣ�k�(�Qf�$H�Uw�	��MiZtc1Nǟ�.���l���? 1�fnbV��,0�; �r�y)C������2|~�������ɴ��%;,P6�+�n�cD��ѨSl{���l��KGT��ս#���TD��#�l��Q�B|�4&�\��>-���/Kb ��tEۈb�-��m�X� ����>����o	?��6�ڎ�kO�0������V�M�
��TD���mm���O��Sd,M��{E>O�#��Ꞁ߈�����9$H�wT�A@�L��MRs���Wa���R�g��8�ӣ����?5��s�x��;�cᡎ>[Uf���/��=;H�g�Dy�%���'L��
�>0Z'���y��<M3[��b��0>!�4�,ѴT�d;��Gq�B{�58�n���[?����q��W������ѧ@�_bm�z����W�=���7_ �Ah���h#g>�%�	9���س�"g%yL������@��Z3b4<=L�����w��A$�%A�l>$���S�췏�d��4��~ �� \G�<���sA����|�d0�Ǹ�����+7*��{]d�6���M��m�5`*����r��D{�.V~E��&�u�rrm��6�F6��Z�]պ`�g\;u+^Z�X
�^;����Q����D�/m1�ᐷP��P�n����H�B�A<�q)x��޲�9A�8��Fpz�8$��r�Si1)��7�/@�q�ʪ�d��0��=�u�j�ֵ��^8q�ȡ�l�q�7�		�(w�n�p��{�'���]c�ϔl)"�5�l�q�o#3��.d���[��|�9W]��&Rr��(P��;�p�����h?�8��xs��O֥e���,�Eq� ����+6z����T#[B���j��� �[L�O^c�<�m�+�I�Q\Y�W%����ž��!��}�Q�Z�p�q�q���]*���z.Ǌ��o�;Hi�����E+��%KW䞠��#U�5tE���]�	�1�������� �8�[��r˒��I�	j{�mp����sE��b>��i��a���Rj�<�˷�C?8�jq����6�It;HB;B�r���[C���q��ˎ��	>���Y!9���+2ǄQQ̷νl��YSF)���h'��!���ӐQ����2>��|L��R'�T��r�.MF;�7̨p��sY	����Ǝ�d�^�Gd�J8�� �$GC����-y����)��>�P�����
F3D��l��%u����.YjkQ	��S��5�
T����}�.���b���Nb_<KQ>���>�,3SDm�w�zkYA��@|�r(4�4�!�V����P�Y�;g��^'�D���W��}~�2�,� -��\{�[���7�<ɠDa�gр<�� �U���3��-����G꺂��Y@��p� o-�88T��0��j"�m'��ڏ�D��"�Q����˳�H����S��6��@���)�+e'`�+ѩa�ѷtN����Lr8)�Q�-��{-XQ�y����'w-�S��S�5V!�η'�v��a��<Ǫ?�?QgFT�NҖb�5���n[L�d��^3��8Q�=���*iF��̭͒#�I@g�{��ZayZO���0/c�2��o���Y|��~Ք%ҕ1�(��,�5��<La�� Z�W�l&��˓�m'���dcw�o
��5�a�$��Nl��P��G���\�N��K^n���k�*��?9�'�z�.�F���2!j��O��zk�۾��Q`@_H�����v�?��::��Ŭ0w<}ނ���B��p�V
@ 5�P9(�xhv�iO�Ex��)��˞@�3������\ur(�*�����;Md�A���Mހ6p�\T�w�)�7��,{�_Y�j�'��v`5�I�2��?���jד�Bx<��K7)S%G��s�&�;Z�$X��ß���śv|��!�� �a���GP�"�9yD��}=*�7fk�d���! �m��O�5q��l�Cb�u�e��=��~��g¾BWTt��D�d���X��z��Y|���ĸ�4��R9H�d7�@�m��<$x��'�mTO��D�ͦ/��?��OO�_�,�-����I�]Lw#۽��uE�����j�>
�̌�^��ϹV��/�ǯ��g_���N!��ߧUw��h�)�(,����`�\&���K��*/2���ZG:'F%E���³b����3�	vBh��7��:S���E�m�<Z�1�v���x��ʅ.H�
��n�
\����k�&�%��O416�B+���EUkW	W�^����]�AU�x��ڮm�Mo�8�O��zn!x�۹��Ry��;�������5��>�J����=��E{U�t�c�R'B� ev+y|���ER
s>�V����c�(�C@���w�xo��49��=�t<��hv	����./:�@QD<���)��G�퍡����(�g74Qϳ`M��j�.�ҫN�[���9;�Ua� �$�4�$��O1�DhbF{�����݁�B{��3�%�=�y�UE<�.�˪uO�T�ZS�]��O`��f>��'��
�o�=��W�ý�+i�0��
�tn���+��p
���Bkn�j���N����x�8���pc�5+��ҵmw�p<�mm�Ù*�qA������v����	�v�P�s�/�T�as.����x����ۜ��W����ׂҭe�h�A�V+���U�	_� Ӗk_-*O�OwJ�P��X����I�\�H�$8�)�S�N��r�j��d9�Z�d�%����@�rH��VEj2��r���}b��e\��`bO:{�稰�v�v0P�d�̬�p��	/R���C��22�8��5���P�У+���NU��`9��-d��ZMB��ΑؿC��l4��,J���C;�Ķ묘:ީK�������t���d���{eĉ�5Y^�<�e\Z���*���#O��Xu�$�q_c̵1j/��	�`�d~�T(MA��;�����$�9��h����o�d0��Rs�=��5�*���'�Hb�Lz!5@ %b�����_��k?�8����%G�X�^.O35��X�AFr)�	o�}�/S=�m�y'L:��ۖ9���/�`���+����"�1L�Åj;XWe\�Fu��j��'
�H�)K)��O�AZ�*�� ���Xv���`v�#�v����y�,�3��T�"�~9W>a�I�|1y.K�3f�^A�%���)�*�wU�|^����|tKS�����gK>�ùzQ�l'�n�'I��L���>�{�0\}�]�����g�VG�%��;�W�.TGy�vO �A9��o_h��x9� �DL����h��mnJH5��]�&�<�k������]��N��P��V#{{�w%0�8����GB��FM��	B������2H�����X�etz��ޑ������x,"���q��%11wh�Z1��z+1V��� ��� X��� O�2T���OJ�����Cue,.Q_�Ր��FS=�'��;�Ū~��� ��щ߽>�?o$���<�� �S¥�5}��d�H��.�I�;M|w�f�V�hL�-Zc-��'g��Ҧ�Z�p��f�!t�;�%6x75�b�Gn#2��}��>���Ѵ࿠NI��ځ����&�+n��S!Y�y@�������LZ��$��M�����i(�W�|�c#�(�l�r�ʑ����JjV��xDd�lޯqEqL��R��MR�~56�j?p�bս&��MA��l�������P���px9S���`]/0�w��G6�]�y?���{�s�	�DnFek���>��RP('ů�?-BTE���S����Q��˳�:��R���md�@=���,�Ț���,��V�Q��1��!���x��N�����v�R�Z��|��MBJ"/�驭.��cU���X���F��瓐�Ң���lI��y|��B���H��5T;Ջ�:[�l�2R��Y���?���˽l
�Z���b.Mi��wS/?�Ж�-�˹�Q:��S�C ��y׾GQ%$�jz�P~F��&U(s�x�o�=��k�#�����Q/
ם���`*�r�-,� kɠ� N�P|ʌ)ҥ�=fdF�g��c���/LMS�Y�������8s�|�Z����0T�E2Cvg*�Ϣ�mmƁ��wrt�Աٿ���:�[`�d/����#j�<��`&�pFB��HQ�d�����w�gm��P�-[����6�t7����J�$�|(�"�����")�0�����rA���)z�z6!��k� �{O��Օ{���𜚥U'������v���&�	��Z��'����[�ꓙ��¶�[�(�n�"�G��;�i�P�d�D�%��c#���vv��]Sy��w��*�-t�~4T6���#�ѧ?&Є<8�Z�����L|ws�jQ�s��w?�v�f���o�_}���o�BótW��{�p��Q}v���'��2����7-��줱k�g2P;,&��B_Ϋ�_v�AH�I�I���l���^�Q���v��u9��mŊPA{��0�L�0n@�魯#p֜#�����C2��~��������衆1ƭcEtثx�A��cV&�K���>i��d�*���(��Dh����ׯ���i+��l��T���%��ʸC��r��On�v\9`�[W���bW������&�#�����[��o�	�����׫��s��ؖط�G���g���z��b��7$
)�m�H)%�W��燞��뱈_D������!t�������|�`i��V�#O����*������j9ϣ�g'�3�.�]h�\���a�$4<!KJ�0p�=`M��9�<������:�k����@�ૂ�9�m��0+��3M"7e�s�G�ah��`���Iϧ.\ٸ�qMh��A��_��՜�a�	~�ׯ�Dת�cJ��H0n�c���"dX�FC����}|S��@L!Iϩ	=i��t�l44���Í�z�b�s��+L��G���9���S�x�s%@���H�� �\�x5_Ub�
5�˴��u���0v;YV�G���o��M���@�eU��q�(.uuZ�{gU�Mή�셕�.xXGF�b���Y��E��6H�����#��R&�^�Ϩ��%f����He�z:�"/��î����ۖȋC5����dDVX�*Յz��hD�gj�-�k2�-��[ޜP����&G���ŷ��X(�?�f���K,�s��Dź'n��#�{:�/��b�ڵlL����hJ�uV
h̴7��WV���~(AdlxH2�>�<w�?P���f�T������^cj�c����3+���w�YYRp�H��Q3���!A�����"wLFU���Cn8�h+D�^��ך�:2q����wY�Z$�)$},��.���,wX�
0Ɛ-��|^iu�Ymē�����'#�eJ���#��iZ�4sD�ڗ�A"�6m�~o�by��VO���N�vB��wu��0�ڼ�h��tT�GD�MC�����r�I/pɨ�o�	�i�B�(m���lqK�jB�R��YєZ
76U!����ñ��M޼Cף�� �DwP6�Ë���l1zq���m�k�[�Xv�E��Ꞷ�����ݽ-Dy7�Z����_'�%��>�6�9k�/P̒��~g$��KUV���l��������4�y3�(@;}KBY�b�;b�Y@HAʘ��	{CxX=���lp��)}���ɉ��n��n,bϽ�!�Sr��5>���Sq��UDX���0�Z�:�Uz<�4�e���Uw@�R���T�N�i�-<[W�08(���p��8�$j�<穀-j�}چN��-=��҄5fX�+��S"	�8s>xj��m�
Er����_����+�jr{�:��y��=?�ӎ�T(��}C��+��
�:*�M%�ܥ�/�Ժ��5\�*D�D�7Va��AZ�O_��w�]�=&!<de��
��U׵�3���
36�@W�ˊ7k��"����)=.P)����>S�K�%���.�ե��x
�5V�ݞRI6�C!��rdb�\�ԇ�H!QW[�3�?fx}��:Xp�-��@۽�e!ڵ�Y"����Rc����!M*y)I��q%�#m��~�Vֆ��,�^�1�M+	EjY�+�(4�&$<�\z�G�����4��� �����-<�i�'�!q�A�Є�O������V��(��{�)�9�%N��v'�ϋ2Me���h�J�}$g����������D�TL@+\�\��S�Q�	y��-`L��Vi��Bp�.�=�S���0E���@71s��E��9����2AFX��;���5r�f����~\H���M�*����oQ3~�������4f~�e�}+�g3b7=m�7��j3�b����qdO /TK��ؓ1b۵'x��r,�~_2O73��V��fJ�{I=��ZQ��z!��H�[�R���|�>8%��w?�c���"b�&*������(�g+E8���`���X�)S,\�V��w��y�:R8��J�2r&�Vb�@{v[�H�;��U�mh�"]�|�r��?��.�@ĩ����)������1~S�c|�Q,×�˱٥��9���G�$ Ȯ��ֳ*���v^�D�6u1�̮((�|��L�KUTD˗0%"����]�u�3��;�EI�g
�"�y_~v2B�4�;���w�|Y}.������k��mгu��o�$���r�·�ͅ�Ȫ�D̮�-����R�v�-d��)M�E9�+�)�\�BU�$���p��i��J$��@"���<:�G�RU������"�(��K���YZ�փJ�k6G��	G�2~��:�`�W��Ս�O�ٯ,'O*��4���S�!e���@�z�ر��4�n���>���	�r#Nc6�FJ�\�*������9��R.ӳ�&�Jȋ�Tup�Ͼ@�1�ͪ>'Tf���W�=`�x$|�8I��]�v��}��1��&m6췁��;_�fr��[?L �ȷ]�	�B�"�Gӓ4#j_��?�#�"_>,��P�,���@�*�|I�F��
B��9k �%e�M��հ�@��#�����d�0���s6r�ك�D9��趟�kv�����R%]�kV/,�l��:��w����z����xIr*�#^�{�ea��@x�������лs�5y6Ax�x4���Ru $HWA����Ø�ܰX?�o�k ���$�E���t"7�%��ԋ��:n*��.&mҢ�W�CI1���8}���~(���2�`�?+Z*{�f�͸���n4��I}i.��ll/�x�Q�G�#�
�[M�h7�ѿ���]CZ\��Z5�	.ɰǾЮ�Ą/�qn�~�4.푩�{FX�P=��Hx_�'T�����:���l����A8��җg��3E���%c���w=SO�>hM_۴@�[M��k����3�:J�{�f� &�,�_�����m�:�F^GW1>lo-�bA���k���4Abr�2��&�k7ƴ~Z��r���~ւ]���q���M��H��0~3�Wǘ�.�r���{~Á?�n���Z����>���O�%�W�5*C&l� c<53і�o���=a�M�Q� CL�`d9�l��H�U`H��fC��g=������m�=&z���r2�dk�R^���||1&����{�f���3��Mp���h����
�b�7
�� $'r6�b�4�F���N���2j�b!�w�eR�̂&�{'��s��i�K�����Gn�}�_�G2Wig�2R�V�H��~D��Ñby���/Q�7�����o'i�Z�R�� �vz=�ȶ��EM'*݀ ��W��R�C�npV�m�ncɀNt]��{�.,�^*�%�S�a�[i+!\���t=��h�����'�=0X�>ZzW˷��9�l�D5W�'�:�.,��Fp��AAa��c-�Ogy�M�_N���Z8��#��M�<0�ϾG��Ը�Zk*.�Z��WߞN]|�7܍ˍ�g�p׃[\�.6ϛ|7=������{�^��
.�y��QB��� �?�٪�+��'Ң���R�  ��d��#n\d�� p;W��ȁf-�(Y_�a���4_�9��
I�3ޟv$�3.ծ6w0���7���'�h��+������7�[%I�p�6�aK7Q��� ����L����QތS�	���u�{�=Të�< �L�Z��u������"܅f_�C%��b�$��l��,�s�Yay6��>�,�W/��GJM�M�v&�X���Cy�_L���I�ß�-��3���u&���-�~>3CT���
���fpk%=�]S@]+Lמ�=�u(��%�ߧ�/�\Lܷ��rP�Ddz�~J��7���{fi��8��dS W�?u� ~ 6����7Q��n�8a���z��^qS0"&�H��o�F�+E�t��}����Gݿi%x�{�
l�̊���iş���Ìu(��"��_�$#�I��Z��O?�(��׭�-��,�S�"�Ch�#@��d�y���� �5�%"Yw�}���S"�����:���ݮ���tF�T��D�&FgO��m�y� ���;	���rR�� ѽF�%�j�-�DIbb]��t�/Z�X��x��E}�x7���[%{d�C�e�mm�H����/.O�%o
)�F�uf	���]]�����<�
�5Aؿ���)��A��J���2Q|K׀����G�)6b��*}���*JF+�ʙYd�&L�ߙ@�;Yc�:K��Q�U����i>�G�������D�Y:�C@#���/�,ԊE�{��������HR����4?�m�i�����oDi���M Q����_?Vnk+*>�a�.N��(�9�����.6Q~NEh���5.Kb�&%��:.�J��"���e6L 
[�Y玣�>G��r��kwo���W:�b��J^�׈�y��9|�"�< �XmHR1 <���H�+������.���#�.I�����Z����f'41>�&y�uu������8���%D`zLX֡컇^x�-K���+�נ����y���=Ǖ3?���2��D�I9���!>Z����Q�/hf��r�U!�骱�I!�k��¤�\�7�7ڳ5l�}�#�5�po6i)�ר6���9��Y�2cX��l"i8*�F�T�x�QŇ\�¯z��b E@�F�/�dċ�J<,p���`0:D	<�qr/-nd�8pA�Yl	ih?x�����b��Ԩ�v�_e�q����5N�C0~țp��Y�B���^9�M�_-���W�3Ƌ\�ā��>~orɈ�7ॠ2��9��g�F����ޡ��27I��tv�}�f�{��s�
��;���P]�5���~ǭ��w;�M9K�/!�!T� B���g�E�@��� �K����Rq�n�á8��+�/��J!x�m�����-���C��x���^Y�����ԗ���3�����<]�l��2���Bm��;{����s'8w%�@]罏^�s�a<b( �獈V�����9��PqB�������	͓�+Ym�BڵBt�e�^<�����s֖��X����:@����X�(�TC�l�Zi*T�vwR9y~�B<i�6~cl�$ή���8�la��$�Ϡ}-�h@!��3a<��D���i�KM4$Ft�G��������v�K��&�h�;�*&�c6)���`���M诇H��/��c��)wo2c��ι�������/6��ϚD��?Y%��<�>m���.��6cK��g�W~�!��2,���$
��0��bk�gـ�~O{�<T�<������x(��sJY3�o�o��B4(����dx)�y;���n$G^� �ŏq��("�k+�K���҅vh�΋���FU�����z���Q�����"_p���t�n�Q�M�A�a�N��D�	�&&�-�Ý�Ϟ\� �[�^��'n"]|R�CJElhꠇL+HC�#(�<��w���b��̟HJ���ۘ+Z�o� ˌ]��>��n��8��#�2�8߫�ν �[���+��~�^��^��޿�i�~��	{�!�b_4�
�'D�#���:Ə�q�iw�i��;@B�ϡ��
m�?��=�'$��y{�C���x�]�^jS�q@C���Y��qM���N�2|G�1����KdVH���W��.�� �4-�p��{�
�ӷzyn��қ �˷�?��G��rD?ʾ��C�NGk�J�d5s>d����]t"G:h��s�3�j�C���V]�Q�����<�'�S��^�4 �7��Z�ǭ~�+S�4Yk������ܧ	����S
ʀ%��x#��J����i��ʄN�����-W�B�8c��@Ol�ݻ�8���+a �2�[�6x�K�sSɚ6��A՛N���oB����i��Y�����~�+����Ŗ��:@,q��}O³��^��*�j\�L�ɦh!���(��@�m�|��k����m`�āLN�?��q=�i�$Q[��
;.?�j��UrԖ�]!7PQ�?��"����H�uEVE+�I���������"_Cֺ���}t�Fo�Q�eY�8[`�3���M�M�N�x�\���=C��C�n ���+=� #�"q����-|G󸙂U�0��Ge�����Ӫ�R��C@x@�S��\PV�����y�,�����G�T��<�
� p)ȕ�oy�u�F&����^k��2����M�M����\p�㗵���?Q,�S{ ��>���u�F��;����t�3�Q�xCLls�侞a���!���JdD����L®�@
X(*���Q����Gv#��K�I��]M���'���7~�����h#��/�0l�s�m��bwX���"���	���zÀjZ�BWj$`w�����F�cW�˿#�I(_R�Ă����Gc|������������@�u��1������`�����"���O͕����~�L�;�-=�� �t#��5�1B��U�F��h0�t�Cu:�{�i�&�|aZ�Q^1����.O�"�tHY��H\W�m����t�NcmOb|�wor�W���Ks,�8��_�uZ�
.mj�9����E�a&�0�R{����$��j���?à:�}���$!� =2��}L���xֱHX���B�.<�ҿ��*e��7q�y- ��ޅ�V`B�����H>��؆�ؔ�J��ʊ����[k	�����	e���;� �U'��9�uDOWE�]:�o�n�B����zMB�Dcz(n��a�g�V�W���܃}��bPk �I�`������fuq��%���^����u}4ß@D˙_��"��~-W	�1��ӜV�vC��-�p�#>|AW&��ي�凶�	��&:[ǘ�u��<�)����L���Y�X���i���������}'x��I3z�������=bEHX�7�8��)	J�n��6�.�G�:(/��=՗]�֧8;��b5z�#+�BM8�QG>�7	F�l;�N(~����w�1������"|r4F����-z�#��m��X��1�3z4��.f�t����q�vd=�
-�;�а��x�T�3>�Y�c97����.*w=8b{q�Z`!�?������r����kR�@N�&��Hf:�Znr�K�[���D}-����!�*a�r�pظb��>D%o�hQ8�Ӊ*#�f1��@Oe�2D���0���XQ�|؜Y,�_���ʍy�9��O���f0�Q��h`�@�v�ǟ��Rm�j�>ڢ�H����4�BQ$U%Ք�p�B7���� y�W���]���0����,�l��c?H	��.!�lg`ӗ��
����2��W޲�#��)�/>�PlD�n:͹�,���4�H�Ӈ"���`?:2���m0�+�a�2���;U��<-��"�D�79th�X�2�w�ZI�aS�.�����'a�S��&���"�=7��M1I��G%-b��J�ҿ���}�s�W�n���c�z"��9$� Z\ �l�^[�����E����y��a5Ĳ�U ��A�>m��Ů�T�O�	{�F@܁?�Y|㑄��^Pg?Mp��� ��~�{	�iu����5h�c����aI�$[�K�_ǐ�"�~�,�� ��)����?�+ �sO��d�����Ѓ�6[���$P�����9$=��{�sp?#j��uK�YX$lFWz�<�KDt�z��e��U9t�xՐ�HH6��$4n7�2T"�f��
U�qg�	7��g���Qg�Ssy��<_�����t�,i,��K��C��#��r�#r_<�w�%���m}?Ҧ-�/[۔ұ���)/���0��̈́���2Ԑ����`x�,��oQ5!X(x�֌B��2�B�W��O��6���J�e;7D�v6v(!qh��1>z!d��NQc\eL��KB�6/J�+��
o��'�LY�m��5k��8�&9JF4����9�Y頿�]c�s)o+�'1h�Aue9Ry<R��3A����A[	�-��W�B��A%/�kеc�\��I'Y��2޺	���z�1#����b��@����1�}����w�6~6����+ �:��3���}4G4s>�uLj�(hs���[6C�`
i_DE,��P*���C���͎6����9~�GJ��!jQ��.qn���g�����V��B���!޾\.t�)zue�tfk��l��ԖI1Թ�=0O�s�/P��)#�4�lmQ�Y?��^�>��a��;ﺪ~���6��/X�q�Y\�nlM���z�z:>\��/G�,	�M�EJ;�����01���J�6�_x�V����x�H�
����#٪�]�P^T^߶е0f�p�ߗs�>�����boy��3W��L>Vg�E*�[.~F�������;O��/�q� �7+j/�+��1\KaB��^Y�HG�������"#��F��Aa\��'K���`�t{��q)��~�k��X���r_m��Y.̴�n�ƻ���CPn	EՍ�1��0H� �x8yLg�@���w�����Xrߎl���^�f��|°Z�v��ȤkS�)!Q$�g�G����0���t^s�[��i3Q�eD�,���7���}���y��?�ݜu���|�_X4��iZ.-���hrj��]�MH�H���"���{�3�SF\�G~;眀����͡���LZ��QN��x2:��L ��1_���U;��e���n)��tP��9�B�~�@mu����t�t�agz�u
��T�Z�=1
>�Ж���Nlm[
��f�)f^�S�U9+ߩ�#"�%K�x�6�֫�9�,EeZ���
]`�)Z5aꀅ�p��\z��f��{<W���n��^ku~�_�Vs�3$j���(�C=�灄��F��eBڔ���������(e����5�!#�9�VějgM�m� L�5C�;�~�����'�ð�
�Ѐ��ɬ9	z���<���:Yd����vTᲃ�	���ˋ��C�B�|�!�����;{f���ӤY1�33�`���w=򽍒�)� ���3��2�@}bS��M_kç�i�oM����⎙��Vu��į��z�f]h]_�W�j3=`M:�_��DCn��C����5܂���(���A�/�~b:@�c�C���e�а/zs���
�$&�8(G�WHZ��r?TR���5�ʳ&�.�.����2(�O��zT+��R�O�ؔ5�]�L�
�c֨�"rSz��j����2�֩n�Pc��B�Gd��[�]E��hnu�L� 4i�d?����di�����X#趬����Z�'�i.�c1�D}����J�yaK�����-/�2��#�����*��S��+S���ba������í%� �ϰ[��-��'�y��t#�F�A��0}Y��w��=۫*c�`��PΟ��[���A[�S!�؂�P�1b���g��nι0cę�>���P��>�jk(�,�����$cܐ����t�Fs�����ޯFN#�K�K'��p�N.��p8�����Z�/q��Y��I�Lb�7�Z*H{Z{^qg1�%ϯ�'�Z�l�;�M�� ������0�=�J4�GKԫ̘���HVRo�P֍
ol�=6���:��υ�i�d�\	�'�r�z0���y��ͩH\܇ dkш��s���A��I#ºv!:�;�	S�
�Β�_F�輯���A}��嵲��u���ppu��9��qoZ��n	[J%'�|�/�m�]'��Ŵ�w[Ж��k�&)���Ab�%�ٵ��Z΅�>H�7�5�d��򍑗P����+�0{^�*U"��vi�U&�I�`Zd�
���������a>���4}G�A��C��Ú�i�t�,:���(�(��֚-1ؽ*@�l���)z1R�[?=�.�/VA�ƣ�l�3_״��V�tpx���=��Ì����7���������Z|f5I�a�4���;Ðl�!��Z����<�&�vAow6om�H���8~JV�
&�A�t�&����[��eb�}x?���+r|������L�ڱF u����c$,��F����݁7F����W|X�n���	~���׆�C�CՖ�x��p�WhPO`���j�8!~J��k��v1^���+�,��r��7����K�J���t�c��[�2vt��CEs�������|٠�Q����a��ښ��d�V6V4�C�b"�,.2�[�'�]̼ �+�CB�}y������+ޢ�E�Ǻ�7=&v$8���9� a��9�n���(w�#���ܱ���{ Lb0P��ފ�%���M2f��R3`�~�<�3��m���g����[�C��P�Z0�O�l#�� E����gڶ% �m����Τ�!��&]�r53�?�<����Jt�L6PּA q1h�W��y9����[G��=}����K�7�������.�Ӈ�<_��G�I��(/�og���'t�ϜGd�_1�W��,Kꮳ��0��,�P���,��S�`�w����n��S)a���_�
���ή�����J�-M�H2������e��}�j�/ȁ�2��:Ý��i�
��W<2�f�C��!�8d~L�2���H�gބ��e��Տ�U�B�>4B(}�+�x�C����R$�t��]����{L@����/���_Z���F�׵�5�+V�+�ې��x޶�2c��0&y��b��D�Y�t}t�~���NKO�2��Y�i�G��)ԉ��P��Tq%����Y��A�k��]��)+W��C�K��Hy�P�5<�O-	��}�W��Q%�@]_�:=P�L �dbg��P��5��R�Д��k�v�6�' �����5(tCH%��ֳ#Y� �����<��1�d!h�G���,�K���5;[�`�C�%��������j�һ�8�_�֯	����^�O}�))o�r�٠g�t�-�,���챞wJ5���W�? V�Ϭk����̑]�O����"Fj�:ǽ(f���EH�+�1z�R����V�&��g+��A{�Ǔi�������h�)Ŷ�C�P��âc0�]hO�Z;F>?z�"(X�dEߝ6��zO{s����	~-����b�F��ĺ
t���R �>2�e��Vi6e�	��v9� �!B%�ޗ�
k8�?l�?/�4��ce��pD��p�S�o���Q2yŐ'�L5�)��~
���AC�%B�������*y�Gu�R	;%X~���W&<�Oޓj�\�	8�5�Ja/JcM5��ct7�,G�!S��lW��0՚�����I<���%9+g߆����p�E�{�,�8:�s�l�5&�^MN"=�߄�W��ژPn t�����	�ʶ�&����OCHD*�TK�9KF[�k��ag�\��|&�e^w�
i~��4@�v��~j_�kQ:�tm�(���^d�_� ӡ��M^A��>U���D����x]�vm��ƭ�P$�6}�Ď<n����$*\�˱Q���T� �����j��|���}�+0ǧZRI;pe��`�r�b�E�}��W��J�v��h����-�`�o�e�s"�Iu��u"g@�5���J�^�M��:i��.}�UВ�Ƀs��qx
�(Ԗ.�>�,���@A?(��d�-��Zڇy����j�J��"@߻#�K��6/�?�|�����|N'�z�v��iZ"���p�: nQ��u�dbI�D�����;�>��@�o�[m@�J�1�`"�a�k�'3��/��Gf+��M����u����1�3�h&n�Is_��;q��&�")�!�*�5�\ �J�!��>Ĺ��'�c˲�s�$��� pټ�D=���-ŉW;�ǭ[S�O�0<��ߛ�l�ܬ��}a�$uݡ5��R���N5�8������W(	s 5?P�z�q?���D)�fn���wv�9���s�n��`��6NM//�s����8��|��@�d��Vm��~L���,|�b(�ȴ�,�<~�fF��%@'��G�>.)�m�q�eT�3P�U�f0U��  I��,�����ɣ@��bR�yH�Gۢ㶻��F;А
���O�[�o�P��O[+�7��`9��[�q>����C=�R����u��W����|;r����R!�;���@����m�v�j�ʥ�����\Բ��o�+�}Ш~#��Dp9$]��L�$�ڽ��Ő�i>�9h��{�T����d�m�5���oA
Q��duC��N�L���&�����
�Ι/��F�������Y�?�, ���f���'�;��Q9�E�[&bNiRMlP@�d*����S���1��w�[N<�o�_̺�F%M�½x�H)���4V����e������mٗ���]C'��n#˱�Y���RT�o{9�A57��e%�0A����n@����I���Y�>�ohƞF�Z������x�8aq�{}��,��I#�8�R6�/rˏ�GM�;�9e���ǔ�et~��L�vY9�����'P��7�ٌ۬�YE%��z
,�H�]3%B�"s޶�*�N�Q��N������$���Z?�G�vP@�41�!N�m���o~3�"�*m$�A��x����5D�~�r�^�4�u�2��P7 �:6[�o�{�϶���f��Ģ�1畃��lk�[�'Z��	z3��)#�vWȩ���W̑-�j�����MF.�0���1$ �G����d��D�C����'���b��q�{ˬ)`�����z��#�`��37�Z�*'��]��|gPoƔ7�s9���(>�a3��4�G!��ݜF̦f���~��*5��ӈƮW{}�4O^���l|9��5�i�+Lh���[�t a����뻓���@�z6ܣxD\�l��g}�l�xa>��-��`��gB.�A�q�J[��ކ٪����Đ\D�`��,��'�wހ�R�9��;9�C�Q'Y�ʟb2S'�փؘ얒�D�#�w�,t���MU�R!�f8@h>��H��dq7o��1ǻ0�Ҷ�Õ�T(4Gx��_c�쭁�a����~	0�8/�;S�}0<'��|�����}Ҽ��S�D����
3,��?�����?�h"�;��MQ�P%��s�!�͂��H̅��%]���_>ͱ�Hh�|�� �?~k�'��^��3�}ڌ�N4�-D��)����w�� �,tL���d6�k��}$�S���D=�m�_�M2�)S�����Z�n��ފ.1����ъKě��:4ݿ\��ʒs�Q}3Lc̒_���"͔�Ң��X՚pA��dA��C)!�
G���ڸQ��j�ri�B��x? �P�ń�r���������i �.����wB��X6��b��7���i��p�Cn]��g�>�s#	�^���	�F�=Q3��c�מ"����g�X����ʳ_�5aAS.d�T�d"�S���w~A��_+�<�뭥�	9�����A|��|0�J��]��p�
�H���X3�2w��/�/gn����fJ��^�~�y�%�A��RHI��#]�6���Er����
�#u��x`3�o�sV�	�tɷ���E����x�ʁ�d2E�$�a���	�2\��ݜ^1x�2�Cu��I�~q���[���`u�-� Ѥ	�2W��ǀ5�������/P��#�����_*���w��K����43mRڰK����Ka���?�F�!u�[����g$RNc�G|�����1ϥ9:��
�EBv{v��ߴD���}�#$��P�p�7�&��{3�Z	`U�|ńG@��(��������S�Ԭ:Q{���K_���8��<P�ƨ�1}��d���6��>g�_��P��)���ep���'��.�:#`�h��0�~c���)��M�
�\3Z	7b�H�8��߸�Օ.�V��nl��8{ibz�ߟj�%��EG^�;NH�KɖR'�%�n�/���ǝ��Y�����Gk�1s@�8G�Z���s��ӌ�V~�n�ew�tl�����cL��x����Ic^���y\���Ph�Ҽ����&"z�tyZr�4� �,��D��EA��39��3��S��իm�U���!����E�����a��e���D&Q&�.k���Jn0܀���<G��	R��0��`{A�p�������R�"�jm�b}��>r����U܋�n��1f�D%��KM�,B�T�{���ޭ�u�����R�n�>mR� �����A����1Z�-:��+��2W�D�O���q,�+����
��Q���H7�,��rVC���e��K�N��u�*�ѧ��#<�����/r�t����䐑�X}�	�Y>��)�;%9�p=x�4�Ċڦ����C(�h��V����b�
MҰ�H�A>�]���cp�9t����:J@�:�M Z�<��[8���J>����2�>d�J	g{�A��8J )L2tK�[	[��3i�@�Q�$>�� guC�!Ý)�O: .�bfU�r��0����������&rx6�e��>�	��"F��T�Q�`;�(K�+YI�؈����"<�1Y���ǒm��?�U� �`^��ߑ׆����Z
��G^����_����YF�2� dr��7�]�@���e���.����s���V�M�F"]���@2M�Ϸ���`��qoB�a��F��õ��� n���%BQ,�����mi��/��pǻiņQtk�d8]Q�|b�㉕�~�jX���u�\ ɉ�E�����(��G��B�)į�H�g�+�<g��?�o���},�71�"(�1ku6�N�
�r�Ƅ,�@�����# /�34sp%Z�L��X�V���tK��4"�R&�i��l�ag���:������8�l�x���l��Ƭ~5\˄xZ_Z]J�J>��%��*5����O&��F�)�w�yҕ�l�]�Y��Yu>�ct`=9(�p1�!�i,�m,�c���~�bu���do�YM���Y��D��^��f���Ay�n�j�2ɟj���b�q%��J]�,2ǎ�P)4�@���3��t��_YA5�u�Qf���K��Wh'����\��W�~����8�x��C�I�=XiLS�y��`՘BB�{Ym+���fP��Ї�=Y�4�6�k0�����Qu�N�2T���}\�oh�)�j:b���`�B5��gy����լ�E�k1Nt���ק�=G�0Nߒ���:�k��3'� Q���®��!>� 5o�[5D熊�}iq<��֭I_��Rֺ�Z���)Ö�-D�E��m��R�C0k&��Rv4���K%N''�&?cr�qs*ja���n)8�y�K�3��Dht�ѭB�]�-�Ώ�Ve��}�ٯ�p ZW��$�P���ZGr����8��g�xj��b$;cR�W9�1NVbLp���~VC������q�ʬ<xgq�6�,�@�.��ԃor�]@�R��]"���D��{�������N��GP�k�X�;^Ё>T���P$�y�������K5�VӐ����%���9�T��B`���ՆU�+A��Iޗr�&���]�t��/�a�:���D�B.��^8o�q<��تB���Ǆ_�?��}�hU�ʝ����I~�T�gҕ!L�U�mڷwY^�"����	�SX�����������gV
L5��b�X3�0Y	�d�Ś@�f����j��>��)3��A"���0�=�̫��n�Ӣ�-�,�fjm���7��Ǟ�,C��}V��(M��� �ٙr����(Xn���04�̼?�L&e`=;w�:.f�-h�~�Q!���p���aT���US�L���<D�lJ������B��uYbq�@��s����N�߰�zW�'k��?y50v�t�f��FS]IJ��Е���~*K�yך��V�7����p��e#��6���)���IU��f-���������bB��*|�7���}�(�dm��5�*���ϊV @����&����!_�J讍�J|�Q8{��qiȊ���V�E6m�[��ؿQ�{d�G���D�}p<c�.�{�Y����0~@l��r����ʝ]  {��0�tFVF��{���]P��Mi�E�J�ۏ9�w���#>s��A��0��g�G�H����w�H%Y��w=p�ٱ�'�a�1�T��T��1��@ �(�4�£rj3e��3�fk��&R$
m�z�*C�qj�E�@��F�oN��s�� T@Ɠ&�n��jhm�q��OJ�H��4̋��;�{V�Q�5�>�������5]@�@��ɬ6׏�SP�A�F.�@9 H��eYZ}�W�2����%������c@��qP�]�kќ���51��բ�@�i���`�����~��_(�؊	�ʨ�:�����8NN��bZ�R,E���p��4k�,�^�P}|hDo�M��7x|�/l�	<�};�0V�peu��U��v��ѧ��������nĪ��s�i-�K�O��r���4J�':�H-���q�?�QlmJhr��W7 ��^0gt�mF�`:)��~�̩o�_�X���jǦ[s(OQ���3���h9�lG)}u�R���H2a�Ά��Y�z��.z�%���i�ʵe	I�g�fPV�A������p��.��!��{�g���gD�.�)�Y�9öcْj:�.[�W�
��LE��q���kY����~L^�]�@xJ��
3���Qھ-�c�٪�&� ]�c������H��<*J.t���|�����2RyI �J/�-ӌX�����]��
Q�e��8MA��S�y.nvĔ����CQ�!f�[5�R��<��mb^�z�2L
TNwO]��������ܷ/6���G��!�JޘK.��D\uY6 ˊ�rwt�:�*Ba�\��-A�YuQ��%mL�wiy	O㊣U�8�U�5�:k4@��0k�[&[��u��E������sI�C1���t�Km��/��y�z� e�u�lQ�Bے�1�lm�*���R����fg>�C�<y�֠���:b��3w���?RG妃e2�,E�:%^�lv�KH����9��c�����q�ڎ�+�̿�8J����!&���r���9�v�q�[E^�����>�|�.��F��%*��F�IQwK�N�ֺ�ߘRᲽ��X��+��Q������b�KǕ��ߢ�JɆ����o~��d��6�>�؟v�;sd�$5���Qk�| ����54����(������֞+�t�]��
�>3E���:��/h�BP�U�n��ƹ,�n�<�����w��p5�n'���� )��N��TsíKr�A�;��[�M���P��Ps7K_�u`�Xj��"a���M����d�]rv�sq�xC52�)�^A�&�o��ԛ��Nb�SY�}S��^�G�ǚ�n�?u�5`� �I�Xr�5����]	,%��c�QxP�T��k�
���5)�-���꿔�!�a�xW�Q��Kk'â�����X	���q�s��U"����ؽ��aWu�7��QHO=�YQ��R��p�����* $G�L�;��5�ֶ+��w��p�F&��)�>ҝ����%@ø~*�i�ĥ�j����q\�n�
��������kYiՙU���<{ȗT3�Կ����i��\A`��F5������%fx~'���5�~'�=~�쇔��_��f�?7�*U�h^���*d��� ��_V�Z)�ϵ��'��= ;�:u z��+�n�+�%����B2"���rq�Qf{FW�@�[�]�Z�XQ��ef��r�|�	��B��G�&�$������X,d��K�����Ǩի<2�IvX����_��*k���6�#����㬋��lj������Q��4�9MQ����1��D����%�(�Ĺ�]AD�e~�,3�K�(�2�V��Nԋ�O,��۫A��XR���JY������׳��a>���e	��������`(���s�!_8��	��L�������fU�iـ�Ip���������bٖE��X����a��kftZ6os��Yo֜���i�:9��M��^�s�7��rf��3��m����s���"P%���(S���kt~q;�z����қ�rSZ��ȁ{���F�
�7��6R�1�cCo���.,�>��m�8�e��^
�ζi�p~�����rhV��B��I�.G���G�ـs��X7 n?u�WHּ��y_w��f��v�3R�P�����i��az6�o���p�Y��R�{w6��2�1����64]@�ł"�I�5B0wbT�����PMK�>)����ET<>�]�.�ݷ����,��ӫnш��M8�s����o����ѺMl�#-��H�XN:Q�I�^��.X�b<�mа��m��(�6"Pϲ���V�(����>����s�"l61d?Y呴R���[1S�	��S�&�#1x5�q�8�3~F� ��@�O�s���Ar�ֆ�>�Q��)��
��}��*4�N�s�2F�����z�I{甖*!�X q�e5�a���<���pj�Z�t-̈́�U����s��[Q'ط��9���4�<��O8ӅJ�P��YN�,�=-N� �;T��s.��Y��� ��@�vrW�f�x��R��!c�l,�%Y`!���[j�Z�6?Ϩ��e�fT9G�l+<#��b��h�C�LF�]�6�@{U�co�7�N���^�|Z~*Ɖ�sl(���{�\r暹�v��A�{+�#P6Pt���5Λ@��*�є1�/����ĵ�Y�875�k�n@m��<��b!���" ��������,����W��ZV�!�3�b�8�A�?��� <&o�Azٙ3}��ۢ� ���ˣ/�7\\��/��x��dM�@Vs�]��|�W��:��P�x�@ؤ�5"c��v�>):�./���3w��:?�7<#�b�Щ*Y���E"���t����]vXj�?3f������Tw��y_����#�HS��&����O�&��PD2-��n<2'����F *	7^2�<��W��.�_���aht7A��t��`�G+<�����k�:]8�l=���#< 46)��Gm3�M�B�o�`�]XH�4�ؓ�=]<�f�ޒ�S���FH�iWo+Џ�Z�g��m�f�'��4�e��?H�İ����b���8/}��_&P�1B~��A�K�_q�b~a�˰h�փ
�Ceu�3��Fe�q� qn��K��ji�*:y�G��Nߗ&����f٨+�P�N�Gtlf�fyK����7�Y�	o���E}���סx �~强 8/ 9���6"6�sy<<������-g4f�P�7�3�7�uW��?S�`�e�~,nYrU$h��"k�Ci<�v^$*캠a�ʬ7v�k�;e90���N�HW~�Z} q�v@�l�.��!&�I�
(<
��������?�O�����{��)���c�M�b���^6�q����+/����s��k�-&)�^���d/��h�����<g��z�3��A3�����Po��Ih��-p �߻��1��H�)v��/�Ъ_�Qq�$gr �X�!������o�%�������[��=��ݯB�vGR�z���U�n�bPr�1K!��1�?���i#T]#�F�ˀ�Y< Mc������65�ǧL��e��i0W�n0��a�@�������yq��6��9�K(X�Cue���zU���{P��ģD����Ƿ�e5�\5\a�w�,T ac�p�*RŔ�P)3�'�ʗ��YLSV�%���9/���.8���U >�P�ט��;ؽ83��FK���?V6u��C��44PZ�I�p�g(2�JG�H(��9�_�3�8SH a����Cq(3$mݾ#���ig@$AZTĴ�l)%ˑW��]�i\�a 7)�fp�'!
z8t���Jz����3�.�j�M��Ռ� 72�r�|���)Z�wU���⃕���"�.ǸNR�`��%;2�������v����z��0#��tS�cCO ������@��.���o?�� ��tAz���M�Cߝe���J�����c:l�:F>�ג!�,�Z1퉬�����g�6�"���(�wO�HW)�t��p_�+z����x�n���@A�¸y���lH�@nB�w�K>5��}�#T14j����g9ݤ/"�*�[�g�0�m��!7U�:�=��!3#���7�O�6ͷ��Y�YSi�b�	خ���;a)�@��R7cg51��O�p"H#��� �_"��F��9OWU�"����cg�I�,�-0�-����Q�0�$+�Cd�,$N��kW2�^��-JI����s��J5��N7q���3w5)0X]�jq��`w�??N����D�B�0m)ǻ��%�)���x�lâ6ε8�)=H����3��;r`zѼ�g�ß*w�)�/`T��򧑰��
��G���T�8�<4r�&��"�(3/�	�	O� 9��.I�P�`���b4���m�v�׎��V�W�z�\%9�n���w�)�=Ȕ�d�'�M�����]$��wZ��*w�z��MI���|զ���P��
.�#F�a]�eT���Q�H����$���{�����O����/����A�^��Cj)��u�[ż�U~�6��y�A'�
Q� �q�����cp`��s�I��c�ӭ᛾��L�;��$�����Y��K�]y>�nL�V��|(J���e[Mg���Ԯ['�	��&�}z�Z��}�br3�&�z{�s^Yb���L����k���P�u�1hJ_RɎ|�ʧ��{��r ����u��*�J�+���% ����H��@+F�U@�:���'�W����k �C�K-���Ţi3�M�n�{�%�Ja�"�ߘh	 +�!���Em�%��&B,�zXܵ���<���Ae\#QT�A�/w��(��A��~�cPK'G�8��3p���~QE��I�z�Y����g���KU�tn<�!)Ĵ.�g&�)��!�ᬮ�[~��9���5��<d���"��x7c�rO�Pz��#�(X�+���1-Cc����fq��v��
,�DO��9w �7U\v�܂іO�<�O��:��NG�%�����4�����8:@29�R9�U��5�,�q7��C���妲VI"��ٽ£��R$��xv[���[qO��x~>'�?Fc��_�1]tQ굏��$z�1����c%��^��zd�ڐ4�89h*u����r��D��ǉ����й�4��ڛYZ�'��L1v��~�'�)�8��U��~���xLԀ,A
#@�A�a���mߞ%�%�1��q�� s#גj�N��le�OJ���\į�e��6`�鴘��N@X��
^fT�H��B@��!��������_Z�C�o��^J���b�[�� ](W(�{�|pņ�+鹶�����*��{hu9����e,�� �l�n�і{�	�r������@���D��ajI�h�p!��fsv��S^���S�R�fe٪�&��j� �P҇<������R���@5���w�[�1�O柂�� ��H�s��
#؄�=��b3N�gITQ8I� �(t�βv?�I�qڏn'��" P^���z�B0��I�;0�d�ET�iN1 �ۈW�����'v<��p������o�ٕk��u�(�@�F�,�v�-�'ʭ�y�tC�Ϯ��N�qi�Ց���f4L#�g�2`<�)�ǰ��|%L@�	;W��|�zW���''>D�M݊>膔���y}e2^�4�kƥ���+x�e��P���5��L���C�Z/�m7"
'}�]Z�N�oFC
���	n�0�c�l�}�lJ��,�
[�a���u�%�`vX36���~���n���a��/�������Ȇ�f����O�ƪ��B���0>�\�q
z/!~ޚ��{�+"�7\O\[���Xg�� ���u�4��fۮs�7�Xv^�+�Z�GT�6��5���hbF�p��X�b[����I��jY�	�0c\�����;��eN0��}���pa+��;��tEބ�(�"��j]�����4.��67.?��~�Y��om������7���r_�[��Dߠ��
d8V��(:��~7�Uz({�{�XDɈNRT�xy�4��f���s[�#�7�u�fD}B����e�~QKvf��D�\}�B�!���81ȭD�w
i����9FM4/���9��‑E�ş5~Եg�g��3 ��Q/�9�U$��9����6P��X{w�iv$]?�->M�[��ǛY@^�"��oT4PM���
�B�z�PH���@3dG����F��f�Mv���ɒ�Z��V�Po�U�RvZ�&�w�C3�9ׯ�>]���|[�*�� �����(c{.�M��8i*܅�c��W�1nK�)��G�k���J�r�A��O��K0ۻ�L�	 '����EH	-BR���.~�3����qt�>B?��]w>
�s�f��_�@�|NwU�/�'�Q�|u�᡼��t���{�k[��F��m����䅚E�׮��n#���m%��T{�ڽԬ{�m�[������)�_� ���Uz��v%��mPv�M� �ao3�~���.h����1��l����q=�aT����O����[�|�sw����+�y�W\v�Q�Lj��xr���a�*�d���,���Et�M8LO0�9�w��[�\ƅ��a �M�+�5�["/��w�{W-K��!G�{+��ȟ�;�ֿo�ZM��N:%!%DS����d�~��zmƻ{t��ߦ��yc(y��N�v�K���)]�uȕ��(��,MI�}P��Ҽ����ߚ6$�-8�S�R�mj�Y؃�k���&J���E��Y�����'6>b��~�C��.�@��B#I~�pp���%��aR��OR�GNvA��$��ع��	x�w���ػ������|�h���B	������'��_�Tb���e��#fc2��ICi��x��._����j��g����?���ː�vN�����o�º4�S�]��>С�p�qW$�����׏*�3���(����A��l���;'�b0�`��Y�<D����%�
-�N���� �|Q�?��rC~ɥ���iFT=�����Z}�UPk닫��q�w��c��3$%u��S�u����U	X��k�|*����m�b´D�"[�~���Vc(:��߁�G�-]1^Y;WPͻ�L:8���$�t:����LwR�ߺ����B5]K��k�~��5�L���� �
hHu��N{w�����P��bs��U �dh��������5�";Lc��=�sa��bYY�n0���z�|~K�|�fڰ�
�V7`h�����ڡa���d3�v�A@���&������ƣ�9�1MD�����Z�qT/O%cw�$-@wx�g�� /����`�L�@�����M� ibU�W~VH2D|����WY�]�=��_0��nU8��>��ND���:2�k��̗�2A��Z4[�+�?�ukN=���o`M8ĥ�_���V܈�k�L�M�C��d,V���V�OY=��J��	}G^�7�z��Z�6E��2Iѡ�^����,�$�������>S�i����a6@!Z�+����-�"����(�. �I�B��s�9|ʯ1��z:��5	�U�%�'~w~/ m?(s�K�f���}�9$Q��4�_��3��vӞ�@���JI�{�߷:��6�lg5�ܞfc|B���A��t!Z*�_tΘn�;e�)��2Qc:��F*e%\B샖c��Sx]�ɮtNT$���3ܯu(����&F2�J��H5ܲ�.�a�X����/�`����2u��.L����Q�Ջl)m����y��'Ό��+���k�1h�b�)Er`"뻫��Fzc�g
+';��z�"��˙h��Y:�(@!�V(j�!7�?�����5*o�<���`ա�����C�������4*p����G�Ю��n_j�-�mWs�yErS����t�bm�����CI^
<i���_#�����s.��Y<01 &�nۧ׃O�f��|b��U�ң�rTKVe�)_%4�Jz#Tz�]��뻂�w��>&t��[Ҩq�S���*���.��QR�B���%�uX�VQ^h$f���yl��˦;��&<K-� S�n��!�/l�?��8-�e��d"��g����_N3���v��=�3$��²�+�yPl�X����a�C�qe���E��x|�NgX��U��҅ �1W*n��%�A��q��m�&^qfn>q�2��������d��g���ސpyK�C���n��x��o��Q;bI��`���{��˱r	�#I�~KK���g��</�s��22�$�C��%��t���D������'����������9�?)~J2���W�g�V����Įk�dǘ�*��7��ן���:X�~�M�W��E�&Ldi���o0��Я#����[�ؾ��0���R� /t��m�4��[����Aϣ(�C�ʑ;�g�w9���d��i��B}�����(6�xw1�������) �|PT�Ώ��/&�r�P@��ˆ��.�f�Z�����njhT�����ӵg����8,�����i���hmk�U�.�+5m�̸�B�[�)�)i؃�j_�$�'�w��E��q8��!����� �:
R�D��o�QȒ7]rKM��f����e���gh,�K�9P_�(����V��Z<���DO�Hq>Xe��� E8��{��Q��8�[�~6&�����Ʒ+��+�-�|~>��87f9���@mY4��פ�ʐz��Qg&�&�a��sN2�E⊢Y�3��W�L���\���� 2dq�&J7�ԉ"�����>`�|�����1��@��4X 2�3�RV$�(Cj6AY]N(�=si�C���J�O]�XP�$��Y�)��%b� ��k�~��ڠ���H�C��}>3���]����~pE�$�1�'Z;%���i���@�-�*������Z��<j��\G;������W�����;�}l(m�*S��g��Y�(�c��}�|	�tq�v�uO�"
�ｅ\�:��F(�p�u7���R�C�b_$r̞��ֆ�ƌ��4}\w�8Hg̅����e����0�_3s�l���;���3:�M���B]�Yj���h�;-ڌ_�^X�&�
sXCk��0�]3������E�A���W(�bf���x�_�f�8���p��F��9?�.H}�~��}��ބ0���h�)Y>H9�>�W!zf�;�l����[��ps��kS~|���R�O��Q,'�D���6����g�� ��ˡs5=J���C�g�]AJ�8�Ǉ>I��T��%��s�q8��N"��jߩ��	��#y+�N�@���ʙ)�����������QE�!�?�P6œ��Th]�sTWU9��;�C*sfY=BD5R�6���ZQ�G6l	�$�;���/�7�VcG3���$;H��n�3T���A'�U����30���Tf����KK7G/I��	�Ѣpa�5�A��M�����:���h����h�7Ѓ�*Ú�HTf�:v<�|K�e*C�$���X�3&Z����Ѯ7�f>|uB�_�3u83Y�*s�}~�m�'s1���:I���зKz���E��*lԽ(�A�o;��h�,���˒oy��?$ͷ���(�=������9�av ��0�I+Ԭ�d�	?�I��_m�)�T�� 8׼׻��-��͈�^��g�?1ʚ��eP�Rk~9 $T�(��s�)��f'�狣�e��� �R/լs>]�q�jP}�J;@�>+��:Ђ ��i"�]Ut���0NE�
F�&[���,['�_C�J�xVBJ��$@�,8�߆���Q�����CEq/h‐gBrXВF��"	cwV�D+\�f|�Q��ʒ�ʞ���c��Ff�4X]��8�(�h`P�5%h~��<Q�߲���ϣX�~������PC&SI�f"�\�38WiN�^���n��q�QV�������D�l���#Z��R���_��� 5Q
[�bA����ĝ���7��N�)<~����y��x�0:�~t��o%s�t
�����+VeO
ѱ9��wY.�N|������ɶ�T~"q
�@ew�ac;���R�Uѕ����̲ƹS5Z�f_�h��Y8��qlw��O�����ȷԋ!:����! �7g)&�eV���4a��do�����yq�	�F����ʍ�5�ntO���fRM����>��7LT/���Un3(8��U0��|�|X�2�H�75H�/���+s�?��U�kO���T��|`���.U�2�-^�vq��k>���G��O�P�ll�܄�@�>RY]7���{�b�/"0��iK-�İ���3}l��[����|n7Ѿ�WH�R��[[Fu�*؋�yWh]�J�||��J���_����a�-$�}G�'6�SV�=�7'��[9���V4`UI�p���nW��b<:[���̓�?,9�����9m]��3���	HiS0�ؖ�E;������ E\٨>���\��p�*�SR���pj"����5�j9���i���__�'FiGL��$�f:X�:��F]p��1�f��'�mX���])7ԂK����裧R�_�	r��p�RJ��9�c��>���w�9���� ΂���ں�Ԫ�	9����;X�yVB�w�|-�^�&1��r��w��)�#���r~��k<:v��v�\DX6��	�GoS���ρ��Ζ� 秓;`>��S{�����ޠ��qe}��Bce4����s��_�Z��a_�K7��׶��֯ ��5�*3/^�E�hI2Z�G��P��^s*˟Xs�߂�������.���^�+`�d��u:^R� ��D�'f���}��e3���2����B$7 ��A�1�H�H��Fέ?�3���B��`�<�o�1{uN*V��&+���r|�gl!M�f���-V�EJ�G��nJ�4H���0���T�xK��w����ʥ�+����'��DcD_
D3�n��xY�3' �.Pa���+���⟫�x~��o�I�6F���%��3}ЧX��@�T��w�V+ �vh�*�e���<��^Jޭrx�p��3G�ꡛ�vs�3��.w\dbh���
�-1 �:��@O��2�s�d�« � ��T�r4:|-��Q>k���n��p!�����g���䃉�P�`%ȬiM�P���J�~�:��>+K.�[��9>=t�c�6wWsp�t���^
JPk�~�ݵ�����"��>���s�$f�h��w�t�+����Gy�_�oQ^e?I�c�R�N9��!�����	4r�0G:�u5<�>�)�]�C1h�5����⫎������՗��!]/"GWX�]���E*\�")�'w�^1�KM!?��ш�Qﯘ��I�摜����*
F�c;##�ژ���̚�@�uߝ��(�щ�&���G�'���L�Ѻ�<�TzȪ�_��Nj��R������3F�A:�c�^�J�	�H�X�ǰ�<�?��]\gN*�8jռ.Ea��E1�-w��i�hX�ma=t%yTt(K'3��c(Q52�^�B�[�D�b;�>Zf�x?p{+S�|6]��$0rn�������6%L��.�#��m8p�0��6�2߃�����*č���Ш�,Z9(�fߚ��L���&��M���aڬ�$��%_ޑG�y˪��\��Fp՞o
��S�%�� �\]]x�`$O��K�J�� hQ�\'
�� tr����9cE�8�4\(�g�;����A�[;�O���[%;����+�YZ�ƌ��4ͺ�O�F ������2�'�%j������F'$���������'���"�ۭ�j0�x�p�dM�,���Oͼl�����_"�H���:2��&�$��:5�P,�,�͔�"Ke��̘��ؔ��"�48`��&��;�RɵBp��M��XB09X����F�k��*�a�h�[���%c�)�����%���F��p��a1�7�c �%���oY
=b�&�I�q��/�DR���f%��F	�RƄ���P�Y���O���~C��놫�����J���y@S�����i#`^�p/�2�"u� �p�
�ʯ���C��,z�����H_Q�?�U'.���e�WcJ8���7���]C�Q$��{ٙ��^fQZT	�>�=��`���z�I )��Ν��ҵX��{���4j�V�~�̧�yg���q2�A{l�]��;t�V�xA	n6h1ӊ.����{�L��j��ڇc�B�?0j>�����ԔS�8�۳8���S q�`�Q@��>�M��x��qF�n_�����լ���	��[g1=����A �Hp>��@׏F��n1�]Q��m��Es-UV�`![�c��Z�`�y2YZ�`vE<�.4epO�?TV�":(֩M=���Y�K����uo�/'�[�tk��62xj��k�0���Hy+��˪���)�.�B��:����N��
�T m�1>WD�.�ǃ�]���M�1&VZ�M�t���h�	�C��Ih�l]6�=bM�� FA:�V1!���$J׬U�ϣD[J�Z{;ʹ'�ۼ�&Z�����MK�">r�N��6yC����Z�rb5��T�V��o@]���/��cFZ+�":����^Nˤ��iNL+�jb�Vf=�7B�G%BWf0�j;�D����T�l�^v�'�_��7N�v��Ոȃre���vYp�+\�kSP-���gs�@�Ȧ?K0�ݾ�JIVш��@�3�Z��l}eo2�1	�o?��R�Wk���@fA\L�^d�\�yD/g�x��>�G鋵���Ud`�r����j���t�ӫ�}�+�/�>�Ԝ�������8��~\R������7��{��n��`SG����׌��R�?�a\K)���?V� Nłq�-ȍ�x&/+������H�x�����|<	�����Z�h ��Ū��#rĨ�{hP�p�����)г.ρ���ҩ��wn���&)ٚ7&�9��`s�r�W7Qe�5���Jm�b�:�L.�`�C��i�u��n'AE.�Ѐ���'u�S�m���	�FA��T�D���ɩTw��N^��TLF�SLh��Lup����~X�t�pP�N������mb����l�����)F�{��}`�8�g41>�'x���z�����\�S48�WK�L�l�̬�a-REt��7H�]�UA=�#o��#]�`s���~���3�
�kq?� weU���L����i��sjtȽ�~�b^�>��DfQgw|1��,m�~�T���x1|P�����HAa�(�ꔝܮF���r"��V[e�%��1���1��,�j�b�)`h�~a�-�4v��e��p"������Ʌ�ae8
�:�0�5a.K��v��(�;�i�1dN�4	�~���lj�\_i�,��h��ￎ2��t|g�\�4Y�@��ȿ�s[~oh�	�]�7 �}�g��jC\�Χ�_��~&������Z���U����zP/��`KWl��y8#������",�Mu�k#,m�W��Z�I���O�^^��>�$��}�F��o�'p�z��"�P��L]����߈�x���8i=6N�}�s��*�W�r���5(��x�`d�RVL�ϒ9N��hUF"��n��L�X���=�*���U��1���ּo ��R9$����nz&�=��bj9�;Ǧ�/y~�B�Nq�-�����Ӏ������ʑ{뭺W^ŧ���$�Z����7�Tʚ�񒤿>ǥ�n��!�\�O���k|�~�D�XmF��
��#0�>Q��>+�H�d� ���B�d?7oƉ>�C�	*�T ��|$J��9U8ވ�J�R��%fJ�K���� ��]���bY4��Kt dpޞ�2X��B���i��'��$� ���w���r�!�Ҡ����nƂ���]��6@��Ҡ��:�8�g�$A�?�4 �#fb�~�Д��!��#�{�����=F���"C*3ӋI�������~��Wc��-x��|ʇ�D��x��d0���?K�${�8�3���H5�C8NF�	�8 ������]uvk���^�%�=ɾ�qc�a��b:��ҏ�9�Ҕ0�?�`���L���̛yn��E��>����#(�9z>�ގu����1Ή׊�W���Ц�
AA]�}��ތ|��F�x�ӄS7�I��૖S��pq����|)�^��lR�Q���O^`5�	�yw�}�7o�K���ZR�MeRHE.�g��Ov!_�$�IՁR�|����"
_P}=���>OL�E�bŉ��3R���n�2~�w�_�bi��ĝ�}���%��U��h	(����A� A;a� e��BR�FB۔U���_�|�D2��h^Ƕֱ��r�޵߸���k��K��B�'d��̐��*6�&��s�d~So�\Wu��'у��a�۵(u��sq��V+��{]�֓��z�J~AL[{����)� ��	�yt�@u=ϻ)�4����+E���4�@7շI�+�G!����z�mHUz=Ce���O�A�~)���Hǳ�S����Eih2�Ycr"��\Ӑ>s���G�m�K]��o'Y����lwXg�0�z��|���>�G�/��{��X�L�$雈٨��x��ڏx�x-v��W��w'���}�w��T"돟�QQuHH�hvV@]]��vi��Y7\r����r�B7����0�~�Ӆ4xh�2�x�λ�O���|�;Z���iUvd�؇��`��H�2��Wj! ѸU�I���Tvl�ŀ��<���r_��<�&���yE�o�'��m~�樸4��<ug+�.`F��B'P�F��v��l������H>���,Z�&N��@@���L�=a�$l)HƵAQ���5x=��JxY����I3;��0�T���&�����M�_Y��v0n�r=z}��D�.)���So˃в"WGSV-���dCP��S�gHץ�]2�yp(I%^�e��)�����s��9�Х�,�@�oo�­��׍ �%