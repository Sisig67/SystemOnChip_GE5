��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����� ����m��Q�D{S���;��ie�9ߧ)������o�A�o:qlQ�����!-�k �|�ʯ�I�gr��A�PmY3t�}��`%^�"��/A@5Yϧ�a?�8��*���p�1/�XSL(����;1fKv���:�N�烋�������}
����~"�ExW�mS�p�$n���MB�X���dLqp�r¤1]��1NO��	���Ǟ�{�����A>���CFĈ���l�TI"I�Hb��Kh�]�����	��Q�����Z�[�j���֯���Mv�Lr Ot��(�R_���,š*Ld(@�v�4���#A��3��S��V3���[��Y"~{�d;(��='R�Ğ�.u�LDV����]��fok�x���琀�C,L9n
�}�q�d&�h�͝T��Ee�^�k��F6 �c?��e���FL��MȤ��iu���
3栍���m��]bM|�(.��yD@�PJv�g�D����ms'F� ,�MӰ��X��Y1� ����X֛�,A�&a=�*��u;��S������$���x�E��0�����v��70��m��H^��\kV��V�v7���i�,M�V#��w߼����g� TLY(��f�@���(���Q��D��m��;��l����B�5�z�L����w��#�����?�z�/$̲`*^�	�si@�q�3�9��y���=I��!A�*iR��Pr�R�.���:�L�͠�$SF��Q��ۯ!��F���u�f���k��݀1�P�(��b��ݘ�y����<�4}��yJ7��s;�n��ɖb��b��jU*y/��k��N|�{{`q�<����zV*� #�C#�˲G�J|ёN�i�vރ;m�W� x��6.p��;P�K�]�k|��k�1f���G�+Ob�������K<s`��t����$���e�8�۪�G��g���Ζ�)G9yZ��i��6Dz��=C"�<T�J6(�gҜKó���F�	[+ҟ��H���5I�m��p8�~���o���^��\ƙ�Su�F[;�x��1��ֻ4}f>��|]�mr~��G��.q���uR�vlŃ�3"O�+4��.��ZWp|[[t�2#�J�U�	9���u�Ê$E�z��;-NU��E����G,u����;�W��������ǬJ\��R��*�蹠���$��>p�6T����G���q�5��1���o
ݛ?�=]c�Ȏ�LL�H��C��vg�s���" He�kp���¥��q�c��w\΁�R�C'V��1����*��s����܉�|�Ijh{��c��O�>���� �r�d�A��[_��K��=Yv��G��	`Zk�Br����e6��O��m3�Ϣ!o[�y�7���k���i5�J�8#�jZ�q	<�����$�i��B���XTQ1��t]���p��O5���gUNJ�=��k����\���_�������x�>����Q�W΋�^,E�&P����㴅�,D��!}IT��C�T�I���q=�k���/�-BϾ]�K�)�`e2�k����|�s�Ѩ����_,�; ^Z���+�T@h��;(�Z�^��&=�B���t�i�a�&b2HV����ye�9Tx��zxE��E�m���1]Ǳh����Ȳ69	��h��W8>��)���;�PN,�`hc&��JVpV�i!�P��s�0����>XRg�����D�6�h˝�O�lor�qa��2"b5��Kl�i���kȫ&D����p�.%��@d�/��У�|S���M�*x3>���o	^7O?�I�\q����S��ᩱ�}���WL��T�e�H�lMb� ��9���R�e�>��p �D���A�}��`�JgW��݋o��q�PM\�ڵ=�b\B=OS�K8yj�f%1
��r�h�;YOQ�o�]��D�U�)�6k&�f��#��F0����寖_һE�Z�r_�{���d��~o����D�B�7;[	]�%C]m���4l)����wA�J���x(��1&�-&�%ϯ��]*1�w��Av��3ԝ��(FI"3�M�<%�ţ���}�L�{T��ib<���Dj�\����>��ػ.��|��a�$�Q�t�6o���q2%.�Q���f���8�侷�2onQ��3أ��H��E�p����� �>x9���P��dt2U2�"�e�6k�����dP��T_�/�#"_��k29�(��6H��;/*��4���e����˺њxq��'w�ζ	��dŲ��p����+~��PY�Q~t��6Yr�"���d�v\�_a�y�,g[��ܰkj��H�Aq��&"Ie�t-؄(+��Qs��dv��x{%�A{�do�'�n�c�G��gp֕,�I2i��[�x	��L����EA��uJ��X� �?�^Ld|D�� �R�RT��'Aut]�%C��*2��t����2�5/��{�eã�9���i��A�R��Vmb�*{Ε��-錚��0�ˣ?��./�� 0i䫢��@/[:||���v3���E\&��8�O���Π�6} E��`PZ
 e~5/'��Sy�U/�C��R�o�6~N2��h)cx0 *g���}~�?s��`=h4�c���uL~���IA�@�yP\*���J��\e&��.A��S���2����th�Z���l;|�BO��)�[3��M�����%sY�Mg�k}�2n��@(��5��V�﷬.��v.��p����S	ӽ������A�WMȞ����+͵�Yk�g�$�J{��KV�:JYxka^>ED��r>��bt�-��1�W.-5� ǜ;US�S-%m,bߍ?KD�ޒ�����~��
\IADժ��+�;��%�y����i�GAc K�Î�TUK�?���ݕ���z+����ܷ����пH��e�Z�"3�}�V�M]�s1����y���M��FO��Q�Ptһ,*ߛYpm�#�S��c�8�R��m�S����p�
��J�w���i�� �ƍR����D�K�>wt@'��e��M�����r>��ޟ���cŪ�zZ�<$�X�I��8��H9�l��{�l�d�3:V��D Y�ڑ8U��v�=��]�,P$^��q�
� Q��:~��2Q��rhN�lL7�����9�5�3^6��{���]�0�~�k=�T���h��_|����?Mr0h��!�GH�ADb�OvxB`]&�/����'��ˣO�bˀD�]T�����t�U���:%[[آϢI�PV�)��#ݻ'i
�]�3p��'o�d
I�V*�+ƕ&c��1s�I���t^�d�oC�}��a�hЬ�X�͂��-�I�7�.ɐ}䌹��j
k���!�������-f��W'�g�dS��¿�3�1��!�t�G�ޱ!��
O�Oq-�1tY#�h���o���+��{�����B������J�'���.���Ї�3!lHf,R�y��p��ނ)"ڻ��w샍��K#�I/���9K�ɵf��,�~m-o�����CWH~�6�*ek���5��������� �J9���'��P�%� ՃOѬ��ׇ�O��<Ar- �D',38�7��նŭ���"NU#_�չ���>��k���Qޓ��
��|�'�t�8��<6a�B<���C��ٔMM#��B~888�5�:���X�LC�9E�yP�5���C��d�Tp�=���fV[��X�`(��C�e��8�K��WtI�>����K�>�9)U���v��x���ѥtvL�*W�h�Dm�z�oOv����h����5��{M{�kH�B�wv���r_�='/�J��e-[6N޺�v�g,��'U�h�.�$J
j�v���>�"��i{L��	mڤ��,x�1Z������7ؐޢ6m�Q��25"M����r��"#�,`H�侢�"��zP��=�Hn��~y�IV#s��>�l�&9D#�m^`����[Z���W�I�)��+�$*� �#Pl�0�E&"?�I�Ŋ��eʚP�Hk�����Ŭp�-���OY\+��;HW��a������J�G&X��I�*!\�Pkf~�Y!Q2��&G ��`����_�iW�煱a ��[���KA��ݕ'@ҷQ�D���I�D�qҡ��I�����-?�
y��y�#�U���E��AV��@k�/��`?�x�uy�>09O���Crg�U<?h������{B�ϣg�؆��E���:�C��S���>�]��v��]?����o�]���8羮��\=��9��_�V	c�~Q&��&'z�tO���F�4��~��{�%��C�吚�8�?cr]�'B���׫���ѧ$wc�//��>�*�����	�3�Iy��wl���u:y�W�\^>2,Q�D�C��K�I�8"�]�_��І��2�ﰔ�Ku59���劗=q�~�De�6q۫��@���J��Q2`ux���\u�Q
��<ժ�̐o���i4�V"]�N�k���Mt�&w8~�7nQ$k�fXE�½x���l����y#��&���3S��Co�y�Y,g�D�s�5l<���L�+ 6Q��=P��3ŧ�,�\K��Ai��x���O���?�#�v�c/�d4Y_�b��*:���M��] ������٧�}�Y��Pm*E<�h��aA��I�ü��˹��+cO�r.c_��>�ek���f��6Hl*(t��Jhf �����򄟆��T[Q 0�O, ����VmIt��qn��o���Qf�@��nrh�i]�Y4�=�%*Tr��|�'��ÌG�h��Ծlp�������a鹧`�xR��C�S_��tS�oB�r���F�N�ߌID�QKwJ��~k��~A�Z�ڴ䟫��"���}�Hx�x%;��?���Rdoo`�˿����D{`�d66�lO߁K��Z�xH�ƄHQ�\�����|s�a��q��"n�
�)�h?�o���Җ��zY�C��(�d���h<�R�r��.ʹ�u������3�(�aj�;Ձ�tG� �͛n�|�T�y �r����c�"yE���+���%���6=�SҤ �������yG��*M�$�Zo�R����'ݟ��W��n��p6�EY�Q�"п�k^]Ao���u�*�2��݁�6[�b,;���+ن��5�?*��-�'8'#�\�u�A��G�b# Sb��X��s���ѹ�؜q�n�Ȕf�dQץC��@���L�H[�٥B�IW6w��A�����n�9�aPcp~���&��B�8�j)����%�l�*�ڎ���ըp���԰�ǱV��W8��F%6=�Vq�1��D����M����L������cfpCy!�W��f�@1�VT�
k�Ū����Y���$�|L�+�12 Tfʸ���G���sQ #��1jN.�ڃ(|Ùh���4�k�;5�1���TG%D�E��s��sp��݈�t�玙(�0	�3�ưP=V1i�TL�)-L����|7��w�oi�d�-�g�P'�	1��}j}��G=�e�hw# �.�w�e6�n���5��f�!�j�k Bo���%Vph?	��E��P6ThrųB�)"�1�w���c�V5��)Y�Fdh���C�������y�p[L�W���������V)�gB����Bk -ES_�՗F��9��T�Y�4xLv�3�z�޴��y�i���)�Mjm�i|O�x	�g'�YzV rL��<�AB��K�J"E^{�?%�7^׀����6(i=fV�������s 	�K���M�ٰԊDͷ��V���^۱�Q�2�[��`ج+gŘ���K~��uTq��ю��p\ky����%���P,ár���ĥ�u��0�|�pg��"s:fw�]�\h�ו�+D��ݳf�<�¾Ӯj��x_
�rI��#1�m�~�ą��.�c��}	��/`���<te��S�p��b��KB\VٝF!q�����;C��|y�8뵞�f�LN~e�b�f�#Y1"�
k�4!����)I�L;&m��UG�w��C&���������7��� |I7Z(�!�� �4Jˣ2I��E�������V�Ht����|$�d���Ag�㹸ڥ7�2�>f<z,�
�G�ܴ)3�����X�{}��ć�纏��ٰ&�$����O�hW��s�恔�+uM/qk:���7�W'{�Þ]�VޮZl�=�:�R���3����,_z����PWP�zV;M*���V67�"O�J��(Y�͵���͈}�S�~�-P]�UcB:�f�m�[�;Ҳ0�6hH��#(�J���Hɤ|��e�U���޲Ѽb���9�|�d��F���Wk��KI�݁R�٤�%78�Ų���7ЭWp�Az�	�.��i�?F�Rs�`�r��j�'�]���3���g8��_g�䡼 �FI�KRL_�*P㜅<���ԫ�Mhjn�}b��!&X����S#?��'w�<��66v�g��ER% ��2��@�@����/��E#�,����}Ln
�H��-��w���悅f,O���%�t�޹�8�֠����;�+B]��5���ﻰ�a'z�<��@���SeI8�zR�U@�O<�b=�h�������!�������j���k���� C9G}( �qf�|��	��*�0�KΞ_�TT˻���dSL���J����Su�O�1�<a���ڣ�J)��|U���#L�Ӫ$�te]���+��&g�	-4�����c��KG���	����j�y|"0P���"���� ��h'�Fپu�8�9���c~�����"̾��2j�N��?$U{JT5������vɴ>�ŷ\�X2��$MbZNi/�}�P�,���J��v�@Go@�ҽ��l/�lYr�MV���>e�'�f�"��q~���i�qt|����QZ�U�� A�m�\4<�)��Iƥ�K�E+�Kf��� ?!�u��������6��rJd�?v翟�S�nA�VM��Ѽ�V�h�0/��E�&7n*�z�Y(�&�$ڬ�OZ�7�"����f�s�|��\
����G�y��Ў2Ā�thԫ\����j)j�œ�P]�pa�O�@	�r%��yq��
��	wT��S/n���w��Q��K�R�s�ĘJ�-p�Ƿ��WM�AaW?�n����'�)?�x�Ng�I�߸���P޹x4FP54^vSĞ/��p��s�R���[��_` �\8�7�aX��Y����95F�[��y���I޳1��PS�i���Su
��/!y���=Kv�.�;�?�Kn�5��.�y�[r|�Mv���>��P���gV3~%��j8-k�"�(�)u~����u�m����^���NY�Y7@��+�M�TiwuK������Ѩ/:����d���vI��Hg����p	?X��0��J�>a�����ă	�M*�S!̓�BVK�p��JL.�?tt�pCZ��CB7G�Zߑ�n����z^>���_�aU$�n8�Q�K�9�tek[JZf��-�,�rfb�m˫��?�B��O�L��v��*C%� *}DZM�ȇ�4Ź��߇�Ug�Y�� �my\O��j����q� ʄ��zk��q�a"K?<��n��6K\�}Qg�^��Y�?r�,��{��e֬*�_��d�W~��;o�������">(N�?B���oX!6����"�e�}�<�V�(�4�T���z��s����:w}JD�5q���!�U9�Ņw�J�;D��	W�b�W #+/���7�P�Z�@U(y�%��fJ�$]V><�������X�җ�3��˂M�@�LO���P��C�@"��'�i�x��:�RbWzg[��[Z)q(̪>��L�R��@�QD@�����ޯ�/�@n�����֎ ��7�jsgE}"^��c�2��(��l�wK�-\ܯ�v�F��{�n�뙆Y��^��L��ղ�	��ϰ���6C�J2 YR�+�IH��jJ@E�Y$F�)���wP&z�!e�Uz|,�"��[��p i�cP��}m��aT�3�N���򥜎U��ވ8E�x9�%�Ib�M���@[�`+lmhC�+?��/���xm�M��r�d>��	e�Dr\�γ�V
���V�e���Z�D)y��6Q�Nq����ͧ��\cw IRy�%��E:�S�p�����@���.�V�;AF��Ӝ�Y�-�`��L� D��j��1>�G0�k�ϭ��&�J�|og}��<f8�l�� |�s��x�<�x
.:@yx����Cc�Qh�pwi iv˒���e`C�zo�>�ζ$��m�I�xk��՜�@�&�J[z�Z��N��9~*�As6��P{����a}�{�Yd��#���V�-����IL����)b���|t2=0�?���-��7�e�z
��_�����F�}T�(�Y�/5@u��Rq�!g֠�x�$��(&W��6P�C�tx|]�i�x�&�1���Ud7�o�%O������>*뤦N�@�_+�w}�EVL�_��3:'����I��� �AʬO�N��V����c즁씛��ۥQì.��#����2�G($Ə	��燃3d� #[n�xX�iEp� T�@Du�e�a�X��G��ߙq�9���D
-�?�X�"5jF�(!���Rk.��MIH�U�
H�%_�ZZ���y�ӻ_]�Kͷ�It/����c��()�,S7����ڽ��7u����-�J,c���،+8P�it�kYcn��=�}�uGMe���pN�SlZ�\R�IQ��������N
����zɜċn<����HJ��۶���(���Jr�lWS[�T��R4�0@Nt�@}���0�r<}Q��/�P�
C+�~��S�����(�C}���X�c����U�_�\"��!̷xe9i���6�#���Wç�ȀXzp���&[��ȀH�����B���	���0���� 50���yk�x4�skBf�\���v�UU$}m;��.3Sk���:�i��y��PA:.��#�<��8�����ǟ��]>7c�
c�m)��e�Z�(k���Uû"��W'[�o�$
S�ό���Tx	,��/�]��/`0����3/�N6_C@�
4�70@���F���Y��@�RGL�\4�W�V[��幏<��Iǰ�ktr���V0�uǡ��(B^(<A1��U�Sމ.���/�Ii4�xX0B��LA��O���qn�Pq�i꜑w3���j�{�O��tsT�,H;�$Y�Ԯ9��6��U&oo��c؜񀽧��x�<uA�D#��a��d���^��|_ d��@�
1_e|�d3
伨��9ʃ2��e��"֓,�,�M� ț4a��K��On��y�-�M��+��}���+|
iw+��'/4�\\����7!N�С�l�i�c:|�l,�l+r'������}�h�������3착ǫ��׀kG��s�!��MY6�g��}�(l��c���
Mӛ�`Ș�u�nl4&���]ĢR���fʘ}�3#̕�K���Z�^||��3+�����3\����x��i��9j	:~�����;O���
��]d��,b�����z�i�n]��B�c�.��T���°1���v��=<[g-��W޴�Z#}��5� ;�Y�H��^	��#�U4.A��1B�0Sl9�m�Ft9��jԣ����=�'�ا��{8�m+��F�����Ӱ�5�@o���4�j�jz��#ᒯE����r��R�}1<���-RF�SBT���ڧ!8��t
w�'<��=� J�)�׬�������,�	RA@�I�0�	s�@@��T&g�h�*Y9�-�͡���"u��Q|&l��'Zz�U�$E� n3Z���Vg�n��a7TWc`�T���N�L<�^�Р�(͜����_���+�'���&?��my/� Q0�J��$�I����$���6�d~�x�[�ǩ�~3y,�G@��u꜈�|��"����B�7�щ�j�d�����nQ<{P{P�:^�����R��X.��%wY��H���K.7T�^j�+Ps-K\i��a���i³@��Z0�2i�~���.p�_��?�+z��.�L�$��:��߉���Q����,|%�3�Ю2<���Pȇɳ7;wQ��a�>�Ck�o���������iV�ph?3����	#�sB��{ZF�:��3lk�QI�ތ"�X�qd$pĠb�b?�Ŋ�CL,O�K�)a~裫(U���#�d_��,���LSazV��H{_�S�nP�Qt���AJ�	qq��I��u�H���A��c�5�u��z�����x�@&�����o�����I'�y4V�Xn��,]�=�TJIڡ�h�O��?K�JK]cD����3�}�>}�%4Kc�a�<c��"���"�g�I��p��y5v�?�(3�.���l����� P{�K��;�O��hE��J�vG��ZQR� ��5�ﻧd2�w�S,)�]�coNpS�Y��P�D}\�Z�ɏ�l`aG���9�Ǧ�ث���T��O�b���	�/exi�ͅ1nP��@Ԯ9+O��I����F����bF@����6g����Ѻ.��3�#`F��+�v}q�h5�8�4O����+U�/�ڤ�B����"�_���S��u�ͩN�f,}�����5��22�C�F��{〼U�R�
|A5�����=*�	@n4�7�P�|d�]��w�lB�w���@K@?6��������tJP��*�~v�z��sK�q҃lz���`�Yc��$b�Q���Ns������e��T�=��UO��qoa�_�j�u�}T�d�:�,�ƒ^��s-�񵑏�>3UN{��ͣUMӽ�nj�K���jf��lׂ$o�~�Xp%a�H���%�[�B2��� ����/�/`(��Z���~��;Cf|֡:	��M�z�N���6�ȺC�lo��g��C�A�l3��ƽK�4��+j�OnN�����#2�@>�9��A��C�ԕ����?�Z8�i���|��L�[g��f�Ꝅ�≈�4�u��)!yu���z��}�	�CAm��y���9��6Z�3�#tY�����f~@ �-���xI�����t�RD�o�Ơ�݊���6$`�G�b,�K|7�O��|�vw민��#��Oh>�ɵ�^M`}C�v3��
)�g�fמ���w�ԬȴYdo:#��=�ק��7��X��q�O���4�\�����l��e��0��+�����<ŧU�޻�ח_g,� �44�Z�U��	���#�ݨ��!8�!r���'AJ���B��<ʛ̕���D�cD	U�BM�B:������?B�)rrC�8�8�b�SYl��^���0�!�x�V.wf5�n{��n�P���)��h_�Va{������#xq����I�ۯM��'��}r\b��ʶh�)4Y,����>��[��%|�'ܓs���~H�$#<yS�L7�8>b�/�Tx��̟�}S��↪�t�SȢ����}��'�1Y�K\�5��s����x��5G�Ε���yx!!��rׂ�	`f�@"O�ƣa�>�,F��n�#݆?���^e��i6>��h���6���mS5�������q!�덌��%�(�S��r-��`R�@��}ʠ)�j����P$�^`i�
x�ݽ{����	�����������L߬�tc�i�zҝ"ʂh'"-y��'�Qp�+I�N~�<������D�4�v������� A#$���W�v������������q��c���Z�>m�#ѐ4�d��2B�}؊Q%�I�7���]$�Æ�oz�/F�T���KM@���%�u�b��C���l�gV!;��R�j�$�k)�k�(��A����V�+��R<��nb�){��Q��R6lxaS�aD�.A��t����bFH�d}�k��s��X4$jpwi+��a�5�*��Ӓ��c/�v�t �!_�t�������
�Y!=�R�����*����������S�,���=��^�h�"�-^	9����,��H���h���eu����zc4l;��ϼ�u^�l���p}^��~f����&�H�r�
A/oS�:1��[ީ蟞�z���r� {����WB�K�P��r�a��,�Ԭ�w��[����r��@�V�ǟ���ڟ
��K�(�|�8X8G@�?�� R@�w�t]Ҏ�Mڔ�w��f!q$1��3�ê�M��"��L{}�}��è���l'��[�q�b����Q�K�_8H$�i�j� }[3M�5������ca&�W�g�����p�B��|d�Tk�ֽ3����D�@��D�@����K�4�I�a�e
T�5��I�qqma�̘]�Dz2�k�Rz�NEG��@���$ь^���N�
�͒��KP�ΤN��=(uP���] �� ����r���UV��<F/��J��60���Īm۰�A�r���9������HV%�8�q���V�ӞvR��k�0|�|S��Hڗ�07�z���3�"�p��BcnF�y�8\�ը"�3��MO��&{F��'��O�3���
*7 ܇�t��:D�:�O]�y~Ԧ�Z7�V���b!�S���}OB0�0���w%��	��MK���S��B=|����d0��O�ő=��#��6U�Ei&��e������[�]�
�ŇAz&T��8y��5@$D��RR��m0������]* ��XF���BR$�����0�k����7^��G�Vѐ��ŻZ��F@�����,�˞Sp`e�qUs���ga��MA�#?�ɂ�H�?x�%��.��Rw�+��Q�O�:��Д/��I�י�+��C_9�|\�]GZ�CW�E��]"$˯^��S��"f��Z��u���>ۂ��x
��5��m����ŞR�?Z����"^)�dU#[W�0`+)��ÌK�U�L^~����c�� �Tz���m��5OGZC��EoctG�u�&C�3�U\���<�
W�����|��#~�>,�zB�3�m[�x���Q��)��T);̧�p�ӏ�P�M�����åUS%/?��kO��%��J2RRa	������TRg4W^\�� �k���j*��Z`ie������q�lu�(��0�vi[�#n/:��!�T��SZ��ۗ3�"p��X�h�W�Z��y�sq��c�\	1�_�p:��^�x���!jK��JGE�<#gQ;���4��<n�-�,!ӡ���I�w�C,�%��#�P��FlX�����$��.~�dmcP�˾l�n�����^��Ah��b �72�}2�|Nz���h4�T˱�L[Ӯh��V �S+L&X�p(������~���G���Y�B��Fb�sP�N�ְ��i�\����.*��2Gv������3ؖ�[�D^f}?���[v�1t�{�st���\�Y|[V͌�9t�������kߟ�K�=��&���q��T��'1h�A�mj��*�l. �vr^��9������X�^��5	��e�\���&U��f�^�Z7�^��̆����ᦦ�ix�bgo<�c��Rv�<Q8�f��Rʳ��mM�Ǟ�J銱+$ �s��8K�'�ΐ&.d�>���`��Ѥ�HqWO���G_����^���~����*@	�_�/���hb�ֲ�u�n:o��.Ts[��R�+
�ۢƌ'%�<Go�%�7��'�qM���E;�h���1�e'�B��� �\MՌ��b)�H��h!�.r_�f���;}�d��k����'�Uk�B��c?�6AbP"%~����|�;��c�Kg�w�sqw=������qο�(ϗ���(��5�;f�ft�D3ă���������`N�I��a�p��N��֘b7�J$v= ��OQ� 	~�[*L	]4�]������ߒA�~��af)5���&�[˱T�ʯ7йse=�ˏk����̥��1��p ܍�aV��:�t�zz+�z�ꑛ��Y�tm����G�Dy��W�"7���P��I���[}����)��@��7z�+g��l�u09�P376��c��]A�\%םj2�U1p���0,�*	@Sr��q��<��7�.�'��Q�Mz�`Z�w�>��w�&�ke�����G��Ő0� �0j5�5L�쒆��?�L�3'��~����$ܒ��KR�����ɖ�8h�l�<l��y�@��&�@��3���ƎCb#M=
G��5*T*��Np�J���@W�K@R����*��� Gud�hž���95��Ϻ:K���Q$��ב���X���7�Z$lkc0w�|�pH�aCt��ʊ�V����E_C��籚�_�H����}F^<�gP��h�M�H�s4:���3`��P ���k��T��^G�v4.C9]�����@_s]ى$����=������������d>덪7�-���_����9~�^�I�{�*�J>�1:�!A<eZ~�=u`���L��$!�vY��:��9R:D�8���,mpF+��o�\���TƼe��\��^�%�G�D�;�/.�>���\d97$�_��a���#��U�o��.�@s]�3��#��~�O�C�102U���(΢�F�[�����|"+�+�Y�=i`K'd� ��q��)�{���%�9E��\��[m�r��fp����?q����m̡ ~e��lk�ƅ����	�0fk#*���Ƣ��yz������B�n��А�J��/1�o�u�W[<ҹt�:{��e�yހ�G����e���	��Wz��V�o�1�����{&��}�mj�'?h��1d	O���FW7�6|�Z���tsύ��,��S���_e�/v�j�����8�|�f�;�<�^S� �a�������v��V,�	��$�?��[2������e*����E�L�cs��0V�sdr���PЌ0aC�ն�ZT��NH�C��X�|�I��W9����3
�h�\���<��Z���[���|�'X���M��p��<q�M]W�����iX �j@��ͦ{Ї.��n���!�����M-ȥ9�\�;ivH�>.�$BX�q�}WP��ڵX;$g%3q�;�9߳�\9"w�?y;o�ga7|l����-v�"�y�z8�(�+G���¹N�/S��:A=YR^b~}�A�����J���#���(ل��!%q�BK�մ��7�l�.+�^�*��ST��s����Fg��/b��w���o�I �w3���v��,o6������;zU�rYV���$�ŏ �>)����6,	h}4ɧ�{;��E�e�yD 	W�=7���tޖ7+��醙�e�}Q��Rg��Ǆ��cYj������%�����/��ˬw��Quش�B�vۃ7��i���|J+����rހ�`�v����8��`C�c����=��x��e���ڪ���ס<�n�l��D5e�&�G������s��L���~O�*A832�X
 YC���j���dS]dm��j:uɠG��Z����c�%�]�EϿ�����	���n	MsB��YÖSyLr�rI��,׋�Uv�}����/ݛa;�|¼��>�����f*h�I��~��J�[������5��Ii坳�S`j�4Ƃ%��h�1cz��|"�#z@��:���i� �#b�q��ي�1�{���%\bq`~b�_�ߌ�d�2�T��@NhP�e݂~y��kk�%G���Al�w3یN0_�<��bR�d��b�0{����]��c�Z5�]�,T��f�n��M� �㑂��m�콊�kF�優9(��TR�`3�w��N��E堁��[+3��p2a��:�ةRR�P���
~���s7�;������O�h���0(�.�f��7���ř�$h�M/�_�M�*��K)�X��ZP&��f  )/,"K/ B5h;�ɰ��0U��<Ma�!r�oxz�M�n�Wj���S�R���1������n;a���z���gY+��~��}EZB��ý�i�r�O���g�r%�.�4�}}����Â���j�qa˱^G�����@17�|CI:��g"~y`KdD��DX�W�!�kH�?#j���GĴ,�c��*邨����� .�'UN��ɽ���	��ߎ=WHl ���W��~~�Y��������,�o�@��DOx6�'��hq�z_!K$���H!����'����¼�kk�F��~
m���z�hW�����I�����IQ���XiM�ώ��{1�K�Ʀ$$y��NQ��&�����p_�
��a�]�X4R��&�;�7{�T�ԝNm*H@K'�M�	ɼ�4�d�pCv�����S�c�4�{�bW8��D�R�P}ާWŐ�Q߃�����&��E�y��Ղ��8�Z5�TR3�h �A�VU��s��1?��G��0X-^��@�B�ދ��q�05�EB�N�ͪ� �G�-4��S�s�(t��@I��Ŕ-.r���`���q�क़1qUMb��y)��Q@�����?�\�L2�������f����2p?B��f�e��hu��pe  A���D9�0L��K�����2!$~�Y�&�`_�P�xnz�AH9�hn]�us����ǃ�[�� �7T���t�Y59c��,ȇ�a��z^,��`|��zpt�j�=�'A(�"l�ahIh������aB��t#��RҎ��ة=�����ͧ�M�qh����c�������oi�ș6�#�`��0N6�V�WR�S8M!ct�Vb����q�T�p�U�ŋ_Z�?��7�t�(q�$a�w�.��ѷ\Bǌ��4����'&��tZ��L]�cĥ��z��wd�<�6�����}�7Q>�M��������Nu"�zr] 3c� 5�<!�.g�S"��}���T#�.��Z�;��/�k��u��9{'�_ŷۜ��f,�-ō-�uS�O2���yJ��*w} .��f �B��V1�3L����f�z���0	F�aR����K���J�E|T(�u�+��d�^4�P�/Ao,s�^�t��x[��+��m���Fx�m�[���;�����H���YQ�9+!�u��l(�󈻃���V��:�t�����^�׼�4	�U��n��y���8=�YMXnFXPGKy��l�n~`�8�c�ǐ�.��%�y6�q�4ߖ�!�#��ؓ�.��Wg^�s�6�VAHfN0�rIl��a�b`�����E���̓`_�{A��~<�>a��-���ٶ^gl�Ħ�ط�-���fF���I�^/��-ҥ3�(��Q�"A����IR�7�mHX1���e�a��߷b{�Ŏ&W�~�(v�-b&�PQ�o��ѫaG3��8�Ԉ����fD��f�T��oZ��uqt?~�D�]�P�Tq���]a��͠�qj�/�=��5�C��ķ$�N+��L�,ҁhMn�+C��'�@v�"��]s{�VX�O�g5����Bx���X	����kB��c�9�H..��g��`O9�遗������u�xU. ;�k���'��/��a�	rU�a�����.�+�<�އ���$6�̾�60/=hR%ˍb�����>j�?ծ�%?Y�,��k��3�Ex������Qd�PR���;�$:�Su�ɇ5�,�pݟ�36�qPF�]8^�gq.���/n� m3�Җ/���j�?Ld'f��N&z;,	!l�q�D�R0��ԝ�_�)'�we�J�����+���W�(��ѹY����]G��9��j5C�ݟIS�i�KTJ�6���?��T $<Ԧ[F|�e`�ً'�����q�ۤ�!,�M.!�1�#;��z?���->r��a��kՏ����sp��2X����ސH���40i���p9G��7�!�NK�Yj��
�t2x�c�Y�Q(�2�	�/.*j���oBn���-p�=>�F�{����>�ޑ|�U]il�	XSzt��1ԃ{5#J�UEȞ���n2��z���M��"N���bp����2�lh�P��Z\t?����cj��9k�Lj^
�8|ck�ҋ�)������?�{vn�m;�Tn(��kڲ�e]��;��3��K*���GT_�����j4������\\��m���b�VDL�Bގ#�(�O����1�^J��k�i>B��������,M�����])��F��㞂�΀��~�@A�d8T���جU}^�TGo�nN@���C��+)���xĕ���b*�%TFB�75���B����8%�{�;8#y�D6�==���\}���Ar�vZDQ1�{�⾂�X<'�\p������>[}��z��eN�`��K/��d�����2Y!1�x;�`z|A�p�H��Z=BA��������E!j��Z�0�Zu+ 2\�o,�:D%Y�\	;�Ʉ\4K���~�A��7��h���m�9�=3����II?�/��K�w�Ů�L)UǬ�BD��>nf�Z�I����.�L#W�bA�eꧨ���P�I0��D���Z��Rq��=�7�ʖ��ݞ�ą�u�lXR��췺LhdO;B��T9X���lUK?Y��z��3��{~%)kF���yKV/�&h_L����	/^?�r]u�mК"�d8�=��u��k�H:ڬ:Zf!
�l�R|00��>u�d�F��PN��ϭ������~�:�7��sVZ�/��la47I��{�9ɀ��	�9����	��ӌR��<;��k�!���k�^6'D��|�,\�w?<��.F��rRH�oE���!����͙�':�.�P�;)�/��!�1��c�hV�+�RJ&���D�q�=�j+�G��~ｧ��;g�݂�#|�'w^%mc���;	�w��T{��^ɞ��J(i哫x\�'z^L\oAT�����ّ(�>�0W��DV �b��[�󩄁��ϐ{G��a񀆴tԍ�4VS�>�S|�fh��MF��4�4�_3��*�'��b�B)w����ٜw t����BZ?��+��*�����f= ��X���cX�#H��9μMh[�y�%ҽ?�Y�#����%�9"�� Xիq�$�,�w�Z�Q�Ǻ�����Q��Jw,��@�
�!w�G���6�������IG�o��EV���O�+���Ą��@8��/�$�39R%�;鄼o�Z���!i��t���h�T/i���qN߇�U�e�yA�͎Q-	K.
��Vӽu��,�+�/�N�1��>�����z{;8_ž��eWp m9߉
�a1�=���dx�~tƛ+�x��@�?���K�T�r��t�
���6��s�I�J���j��y/^�~"Lq7�f\d�����NS�lB	�h����i/i?�O��![@Zܵf~�f�#�?��Q�tj��ԩ#�\���ա�ה����O5.b��"t�BV���':�1�����L/����$��oHT�c�����S�6@�F��dQ��>�LMn��#p��e�ު����PO$�"�;B^)8����U#	�����y`n-8<w=�4�7�)��	<���v�E()n#Q�
tǼ,�"C8b�Ϸ-��G&�L(D��S��_�ۣE�9�<I"2���`��bI����iC�c����9Br#�4�*��I�ڢO�{���_{���/<g���6��S�!R
BV#��e^
C�,l��ט>�1�F-��8m��<|��'[>��NL�|P�c˹P.�J���U�>=��z������\���Ԏ�p�O���N��ΨH�����&�ܲo�*�>o�^�S�a����p�"t�&��a�R�K����8�2�rp�~�����k�lf�50$���|���H�@�nFN%ʮ�w���}��@h��Ԝ$p
�z�o)�;'O�0p�l�r9뽵ۄh�+���J�JӁQ	�)U�tC'��h�X�XK�K�H��9�^��\��#�����2�!5ɢ��S��hM&\��%m���U�V�+G` �6����vtk3<@O,��ן�?�_ x��S���h�F�V���k�A�N"M�{���^#�J$���������"b�Eˑ+BvDE��+K�����3ck��u�1bG���+mO"�\'i�nыz�B�nx3�6��cjs�Zu,��%�n���y�p����]�D�.���?�����HF?��!���W���i��F��)p�8
�XsA<a��]˩�VJ��j���hѣ�E)���[Ď���|,>�*zi���
�;Dߵ�����RF{�[>�Ui[��-�JU^㟄-�?����;9�F������k9����u��d荘���퍝W���K�9)���5�_$i��H��U�^��q`R�?�����ʫ�p��G�d��D�e9�̌A/��t�h�f��Mt��C߬�a!f$_9�G�8�S��]Uw9�
I��сTp:,%�y���R�b�
..ɀ��������E�N�½�ȩ������o�y��eT
��E�򒷨���5�|�'�g��\�����K>�x�����m�����gd�E�\��S�b��<R��H#ǯ�;ot9��wf�EA���h����)5R�)ʼ��w&<o'0E^����(�)�A�C�+2��M�%.q�i��k����O��*�#n_&�,��O��v����dp:�0t)�Du��lDC�\�a���CPUk�y���[QF����"����g�C�B�4g6�$]�\(����aB��4\.���펦��)�~7K ېq��E6�/��jWOW s�k�4|��Tm/K��2�H�)Qo��/���ʘs�m��d�"�>�bԚQ2fu���b�}Y_���T������p�N>�v�)f��M���Pc�	h{�2���7���]1J=1��9'V4j�-���w$�!�����Aɑ]�o �<#��A�5���4������s�h7��r��p	�zPs�]0�� U�N� ?G���j+��՘n��ތw�g�{�j��k�B��[O�KZ�z�]�N=���K
���YIT�S��/�S�?��,(����e�f�B?�fW����׃��Ҿ1Y���5�Լŉ\�mi
�=?��`�=3C�b��gp2UN��15�<&
"�-��a�ᒛ7R͸B4@j�U	��e��*PP�2B��/E�q8�����3T�N�">싋�]D�'*����٪&��I�Px��@��)d(7E:��c^4�^���댫�Gk�#��Z���_�E��nC�]�H�osi kZ�:�X}��ʍ�8�ʢBmN~��4�EĐ�ݠ�n��bY����L��v���9�6�[I\��\��D����F泔�C�Br�ܣ�a�|tw�R@��>�����F�o�:`�����h#�m��4R�����U#�d������%���DI�0�J�>
ʵb�s���C<��Z��Y��|#\V+�ǈ��-�X�5�<����Z�)�*��-�eø�c�G�����TS��qxR��ڜP����/�����M�e�uA���el�)�K��u��l`�h��T�P�iJٮɧ+���0@ǂ�\�)��I��%��CXѝ�Ǔ��{tK������ҽ7�3�}�x���l!=�,��	(3S�F���HS���	�\
|�fU�a��T����%��ZL[�Թ�B�I6�8N���*ů����Vj�Tx���Q������!$���!Ҏ x��y�[���c��
G7<���ă��4gL�tŋJ�4��gL�|��`�C���HhG����<Fm�Ȫ+�x������#�6��N�yV�t5�v��&�Ĺ����_���^d8cV����i�3�[���t]�VD��:Ȓ�!���ɓ����<O�{�S��R��i���+���kt�z%�%��:������ۉl��������n�U$~��fw�t�(S��K?�V���?�eԮ�r�wB� &+jq�.n�qe�j2b+��Mg��nI\s��"8�P���}nq42�K��'��3�=�	B�x/_D4`PYYJA� |�M���	e\�,��I:D���{��DoW�g�'�TƗce���)7��2�_$���]���� �.N������U�j����{t V-o4�(%ZVu�P�$�erq�K=�����*pa�ü���SV^I��HGXB�'������o&ߕ[R�J�(q(HHG�(�|h�/�������+���Z�����{��3ʨJ����z�R�8t���̥ӓgN8���)J.{�zo���o�bs#�޿���]�P�U|�c.w�ᱴ?�lD-��v7M�Y��&��̫Z���V2��p�pOG����O�N�1��Cv"3����"pU�ڴ��)#�46�v71w��:n��c���웽(�5@���-e�ѧ�3x�c�bx�(0�� ]5�Gnc����^10Ԧ�X�j�m�{���]���v�����BX]�2P�A^�l�_�>��L&��]�p�$\Ռ�H_!RcW���*�k������]ŀ�sD2;�鸪���y�6� 
�ؐ6 �Z�9��T�<l����"<)�����M!:�x���#�/��;����)2ۏA{�'�ފ�z�2υ��� ;jn�������4���B'�0Ƃ=�.��|驭�����]�F�q/�g(W� Aw�x�=��/l>wU�>�i�|k'`aiH#��n�b2A�oK@u*l�D�5X�0~X��V��/E+���5��A�>yVE������MN��8���0�{-��^�����UýS���������s�NP啋�ο��IZ�w��W�ٕ{7P�i�a[���\_��<N��#^O�w�j1.I!E_5D�q��R�FΧx�֚ԇ�o�̤��E�.�
��I_m���u�u~XN�0�_��
���?v��8�Q쑅�������'�D��w���;���_G���� �+�w4��i��z����i���j���ЕYɆ��w����h�ܝ�H4������j�K�͙��:�y�ƙ��hIgݦ�+C���w ��ȳS��; BM�~�\�_�9Z����Ş_��*��� ��/�E\�����π����$s���9Z����G��F
9�V�N*ӽ/h��(�)��(�( ���.$_�cґs�?&%��bi$�wv�!��/:�S�v>eG�8umx��L��w8���}�>T�q�k�$���$�]�ڬ�w0�橁��~�>-�P,5��a�0�.ߺ8l��2���E��.�o����7*Ӝ�?=��+ X�Frɐ�ۈ�H^����(D�)� ���r�L��!x�EÅ�f!�>�4�^�!�˟�b����D��v�T�iDߩ�����`6P� ��Nΐ׊$d��N�r;�P�!�D�T���S/D��)	NEյEc�� �R���*�k�w�|�+��ax5鞖�Z�aL��O���#A�6�z5Sz/�|R.	B��%`�@�N����T�/��P�9'��*���l�xZ(�󇈒��sO1�Kun��F��$�zX���?rQy�M�H*g�;�q-`�	�b K�A�:��ae�fNy .�GIk%t��B�L-��)���[#������Ji3�N��A1œ����J�t�#B�G@�5��m7hJN���\���֓�}�j�v��g{UJH�+u�����_�jq�`�ϭQ��a{���!��Cy��΄AY�G�Ӌ�$D���b.���"Ӏ�ۼ��X
��@���,N/f8擉XL�=�M�L�#�x��:(K��ۻ�,m�����f�mĻ'�l�=b������Ѐ��
�����(��������')��L�BT�<��P�2���Xx���d�����?���2!�d
��E�܈�Vn��H�L�SXI �ٔAk�	�|�;"n����ĴC��C��ݑ�w�c��TZ+�S���-�+BB%�D�[cn��$�u�M�1��R�-�9��}�#�H�+��k��z��C�^)c9�Ik5���afցu_\�Y�|����5����F#��;fz٩5��!�{�պ|é'��	�i`�/O�>οK�����A*��Ψ-�T�T��.�:pc�S���A�;�pc�)��`1���{^���4�N�5'�B��� LL��#�+������t�5B�U�-����W`]py�N�o�����M�+�|�����/��"Ϟx���/�r���uip��ME9��\��c�f�Za�~㰶$����9<��|���0z�]̖��9Q0}|D��s�;�jf��A�E��ʘ=����&�Ӗ7�6W�]$1�xi&	��7�����e���	�������ϴ�j�O�k�a��Ɨ�=W3�6 �=�m���a`m�"Z��b���I!���ϱ��d�zD{F&�N�`�
���`�9���~�I�n -���ٕ��=!^$�b�֢iy��Ir�A!PdXL�����!����l��-ư&�h��VX���%y�Z��<'������g�؁Y£�z#��v�x��/̰�����A���B���D��4�C��Zt 7�~����og��݅���z��	��P����Ǩ��Ѥ?�ϔt/����
$�>]ґi�E�1U�<�;^\����7��B2II	]Ni�
a�.,��}d��� ��Rn��3}7�;�IO݀�Շ1m�T(]��b-M�B��J�1� \B�f�6��y�=�_De�����~#�-@K�ا'�FQ<9�eH�G��Z�V^c��3m��(a�
�g^"e̙��5>����$��R�H��Ԥ�z9�\"'�
�~�?7���^y��߶��C@�ݝ�v�X�Φ���|i��5VL/zz[[����U��`����)) �&dR��}.�(���1���h���I�+�H��Piqt����HnQl�'l��\V��^5�W�,�JN�#|�Y��O���H��>���3j���m&t���!���`R���SB3hx�J�!o��W����wnh����Ds��q~bEb�)�S�ᶅ�K������΂��1}亾2��^��%N@�MF1�O�_^�qˉ2��e�J(��Q�F���_����d��n����1$���WfR�$�cz9�(`Ω3�a�H����6����4p���N�w�����U4���S��=lJ1
U��@�>�?��.�1�θӓH��5ۄ ��M̓�7"ol��c��2ʵ��	�a��#�M.�,�E:��<�4���'�c"sx�+ܫ���o[��>폳]3��s�HT�t�J�}WTT�|��t�-J&�	N��qn�<� )��ȗ���'9�n	���#>��
u���͊VPP�6%
�*�JUO]���v��'��-S۲�3hC���R0ϕG^��n�"o�Q����H�]^5>��Ȝ�US`w����K��R�>K$�FG`�lr��'�9�Gc� *��64�g1�c*aMn<���I_��B�_��{�jVI��et��$�M&�����njfÆ�%@�������=�7���h����L /��m�Y?��]}5)�q�*ހs5m���}��٣��U�,���;$Ĺ {��"?��?"�^���b��׍v.߁g"���@���U�f� Z���R��3�C��I]�+.ajBo�5㣀�JS/��m�U;��)�� ���C��ʸ�e����y�='-Y����ѡE��xy���	�G�nۗo�����}AT�~����9��p�"�l`�b�r;h�	��.uW-pg�/N�Az�mxxsg��W��x���b (K�s	������'ץN����wf쑕vq�G�����#�ؐnC��5�j����.�-�E�!g%;�Dڒ{,Ҕ�̚oS��@�~�ɳV|�b� 7���%OqD���ޮa���7Y��&��M�_�`����,i�g��sȲ�9U=� �XE�Q�wɂ�`,���<��oc�O���K��j� 3/4h�I�W��H�����Y�D��B���ů�}3_5�@�v}Vs޲Y�T/է�ߩ�7AwG�l��2��>W���_��k.s�ҰF!+CNpz-��hRwH���#�j[pnW^�<aB	���/��{7�9�d�?C�vV�瑔��;-������Ўd�l���D	W1�C�A��0x��ub�(�"I��9�����O%�EY/�t��,܋]�J)� 6f�00	�/���}mܤ���y.��d�� �zv)�q!�t��a�͛�����O��
c��ߎtG�� f�@ި:%�t��`�����4!X�;H�sv|���Y��Zg���&W�Z��r�`n�ݤ蜯���!d%Y=:N'k�0�mS��Ue �C��0��}��M巨i ��D��u�� ��P2oR���:~tF5
5��!/��bF��V�����VK{�����#r���G��|��L,��Y�EqؒFE��9^j�5�=� `������H�y&�1�]���]�}2�7m��JB�{q-Cu�އN�xA�S��D�A�)�N����5o.}s�C8�u�;5���t$<4Ș�`���������mg�G�dJ�=q�s6=h|2+��Q��$�1p����~:W��a3�����ܮ�?��d�onH3�4'�f�[��9)�%�������	�;�t[$௳F>C�����n#���Q�W"��a�lH��a|�aI6�Y� з��(��x���Y �P���ɥC�o;m�`ntK�g�Z���7��Y� �1��^H�q"w����\G�?ɵ��}�R��?��Vwd����</y�+E�ڔ��P6~��͖����(�΢e���I? w5L���WF`��:Ф�;��*'���w�l�`PO�,�c��+ף4�{
���y�����b�O�s�&��/*V�~�Bqaj�1�C����c%�0hr�7��������G�B����cF_�� W��,�R5c˝�SQ�찲&��mV�%?�y�5�Ѧs������<>��ᗒzn��O����ɥI�hB����&��WS��I��@y_eIaN.Ȣ�O%�f��b㧼������P�,�2�����*� C���ԩ�V�y�~����:�g+����U>;o�34b��p�w��H͞0w���h?�k�'�5���
	��bS��:�Ը�^�	O�����"z1�H���tAh��@�𺊮8����+Clz����F��-�!�6_�4���Z��D5��A�9:�JvdXK�3�����;�0B��5p���4��\ߟ�֋�F[v@��"��4��**'������gx�?`C�q�\��� �!x�t�J�ϮS#��d�� �qS�d�Z{߂�c���"(f'ĳ��
�^>�fơ&5���4z ����V����C��ڀ>�*O�7�����s-�j�d��I�T��z/&�7�ouЮgb�&`@*�(�2Z;�&���]�a�m_��ͼ='������Sa���fR��7�mTXO�
%�U�G�5B��(	[�d�@�s��ԎU�x f���D�J�QW��%��QN����Xׂގ_fn���|�-����keh����1^]1XCq�9Br
�2��O�O��,<�)CK����$`��R3�)�	��.������&ys﵅=�ס���MK��#|͓tɣyih��E�һ���~K$Hd<�)�P$�T�)�y�9�B��X$���L�{���C��bI��܊+�9��|2ɩ+G>
�;�3��y����-J��	�
f}ש�	}��T���r�]�#mi����D{�����Ko����v���<\�d���6�.KLO�$��* 
P�� r�n�ⴌ�����J��'`U]��z~sh����BB53Y�]S�}E* �g��ˑo�Y�+�����K���C����]ҽ����� tC7�`��y ��5���J>uÊE���E��Γ2&�Va���DSk�;٥�������*[�V�(x2�?+`ȗ�R���O��U���4� kD����d�U��*�7�?�- ���b���Y]v0�Py>�`g�m�1����("j�T�Ǉr�u�n܆��q�[��u;*7�Cp(��o@�=�t����ڕep��<�ϻ��]�K�L��P� f <�K�<<<�]�(PW.��q�P$�29��"���b�K�<,�l��|Sp������r��J�<�R� �h���ğ�<�5PQ�Ŏh&=���	�1����>5^c�N~�E��f�v7?r�Rߵ�����
�K� p�����֜��������+�I.[�O3O��������fk/ΐ��zػÒ�(�y۱�إ��_9�Jz��8�oE�{W�ZZV���SxH"���:���,S�.!o�E��0����}4�;�:<J0L�B�X�2�E����w�u]��-s)��Z�4�) ��N�+�$Șy�I?�x9����Q�Ƅ�0�N:��L<#+���+�p��/�������޺�;0�n=�U�W���:}[� ޵�.��ar�5�d:�0C%0hۺce|�Ww�b��h<�ʭM�y�r������E�"� OSJn5��������{����!�u}$���\ަ�ᗑR���-����2��t����gJ��eN�?�Ik�x�?�%x���q� �v��!�����[��#.�{I��,>1SH�?eM(����ߝ���X��p���?�d���j��ܫ�=��XB�$��fZ�xs'�����[���1��Zp� �5(��{�݋��E�$�X�mt?�W/�>߁�F�f�,���<jC��H�u��*ud.��n��T+�t�b#:�/���n�!�Ŀ �^��I�U�ޱ���4s��:�M��I�>��j�t���u�Ŵ�ʧ�<=���WP�|��߈8���	g�P.]Ϣ����N��������H�~,��t�����g����}n�k8|�^����c���6�F�W�ȵ?g���=��f�M-�k�J�����V(���~奒�%��?5{=�3oynaf���@`^���$�|��Oj���[/i�U���� SB�+I��������_����'x��d�$�U��	y�%;����J�ws7����W�
�ܖ$��Z�
����Є�a}s ��^mO�8�PE-��ըe!��(�B���͝��f�,�R�S�e���J+��n�/`�6��3���z"4_4�+GP�ӤԂ�|�^3���a�Y,cd��h'�����u�dtB���/T�{z+�[=8IYt?`�-�:���d��q��/觴�F���q�x�8���6oV�cff���"��m_Cg��m`�if�)�M��C�Ő[�2(���I�H���8�B[��jv��L]83�!�5���P�^­N�0. ���6<͓� r����\w�^�s9����մ%�~D�ɠ��7�]�<�� W��MX�˝ѐ���o4��;����Y9���Yc/�D�e����بǈ�����O�A���h�8Y��_�E<��[5�i��wE$�ͮ>S���D�a(��E���|�h�KXo�S��;&WAK��Y׳�Ն4P3��XIl>^�!��j-C���xM4fU�( �R���v[�H2*ob�k�MΆOpE�:�
��"�4�b��l�����mc��K"����������!C�r������؍E��p��~�� L��E|�҃�S�r!����In��G�Ѷ��8�qc˅T����\)�2�Ƒ�f\A��J�t��A��0t��z*�n�p8�U�X^�.d' I�g�"���T7_W�j�YRh��?�U0�qG��zW������9���I� ���ڕq�� �T��Xw����K~[C�|"��D\�^��d�:����䬸�ަG�X�ѢO�FP�=6N�e����U*P2��y��ģ����(v��#�8������ޏ�(�+X���&�T&Op�@�E�-ꋵ�r	���.Ɋ�oM�#��Zq4uUv='F_��U7] ]n01L�[�Us��[F�m�P���(���$�0sq9�Y���ta 	rwr[l"���K<�*��!ta�*�������O��Z�lr��)���gÙ�>�wK1���U�}�B\���dC�_Z+=��z_1������ſ��L���&CG=)�P��sQ�+�����Ycf$��][��M�`���T����D��lܛ�KOv��X���w���1�p7X�쉲���(d���Szͪu ^�N����y�Z�5�$��Y�����.#̺�?����	��l����k�jƣ�V��)Ŋ�7J���ۨd2�N$a]'���v�iIZ��S�s �J��j�I�hP&Y�����6���c�� �U!ν���PQ�%�'��i���X��Z(uh��
� �I]�W5�H7�^�RVb�{���˹'�̶3�Q�o�΄��xl��c�#!z�E� �G.���P�Q��>�C�~k��-��>Ҏ6����=F�ve���Kx4�1�%^C���%�Nضs�%!��W��I&�����)Ƿ\H�Շ��W7�n��$�	K���j���F�s�|�M�|(�ERoJ;����-�x~E��+H��7x�� ��	�(E?E2���qH�Bm6�	S�z\\�u��4S2���:��7��y�`Z�}}����7I3�$�UA�̣ɸ��n����m#w���d�[�0j����v�̷N�����W\ՌEJU��F�XK�%-\�fpS����6��S��6\�.'r��h���z���1�aZ�#��m���T5�o�6�lgY��ޛ+�997-ֈ����P�?8\V�P��e��s�
�o��H0ž����M� �P��6��%�N�T�w4����4M�y�?%�QJB�a�b���7p�gl��[���.���T���O�m@����]�._���}��s�þMWɺ����=�'q��hMc�E�C���N�G��p?�YV��&e�(IY21T�PM|��.��59i�r��>��b�E��'	'������a�e��O�{ح/)�ϙ����m���<��K1T�%K�Va��M�w�=���7�|A���I~-4�t��r���o!�%�����%�^�<ٸ���Uۅil�x�g2tM,6$H�Dq�`�/7v�B<^^p�r~:��D�O��bFýiSP�Z3UA}cS��r�u���{�;o�q��+m���[7N���o}�;��.쾩?^ɧ%�P?g�j u�r�ی�K���E"Sgz��x��S�A/�0+��)�%��=���=MGAy������N>ējQ>���Z�/%���4�KK�?�a��YP|�]GOb���.Sd�����O9���up�|T|�ͯ���#�6�T��Ҧh�)2�'��O�%�U�2����?C%��c�0�5�������ubSr#�j���*��Q겺�J�2J��@�#`/Q����d�
6��le>`���O(Em�VD�m!�⬆�#���<�0X"��h�ކTl�$8��)T�R�����l��Y���v���Տh.�����F��0����Ϳ5��M��z�azu�Cr��(V�zFU�Q��������V����ű�e,fq��F�-�f��4�cG��Si� =`�ώ��$�c6�_�fgc% s�aV3��3ؽ���:�`z�b��}���L���9{�����P`�zk'��l� �2�!�u�����
8���L؍�v���W����8Ja�s4o�HM�{���I��+�^�gi�s�\�� ��;�ʸ�l�1�2S�W���px]��mϧ��C8	�a���xl���A��y� w�{JA�.��hr�s��5�S΍/aqU�ڴf��i�_��h�8Q�5���F/�(W.�.H�%��Ѥ��@ D�mf����4&VA��ݒ�s�-
z�B6L��qb^/��CE�m�0$��n�:~��K�&ŧ)��I@���ם�~jc�bV6t�_���k2�Z���䐨�댎3��M;�~-��õ�
���3o��t>a�to�}g�I�$l�y�����sG��^B�r*���V�X�Id�g�X�K��{�w�cM�A�������T�YQ��:x��M�Q��e뽉X��m�%��)}�6�t���RS�ɫ��|�$�ۅ����c�`�Ma��]7�!��П	�qۼ�'c����S{~�?oV�m��"�����>3Z���^Mu�d��c�����VFut�"�R*�J�~	��1��X,���^77��J���/��E�M�ֽ��
E��bJN����$S�F����������d�Nȳ��f-!^N����Hi��N�e<l����}[%>�>����6I�d�7��v{�;
�K��'�Ɓ���ٝ�0g��eg7ވDa|P�j[�u�{���ꥀ�F�܊�@F�x/����'e]Y�P�r|�K�77am��C ��p��v s�f�^3n��&����RgP24�y3�UE1.N�a�6��;��"���wъVe�s�d�o�/����[ŭQ�8n�{����0�>�п�����;�y�=�? �����0v����w �O�HbM@�w���$��M�����Z�7`Q�5;+\w���#L�C���qZ��Gh�����N)
[�~����jc�j�����&����ؔ�3X�'�;�8E��%�Ѝ49$�l�l��c*���QJ��>�ga��䰎#UyqiU1�ٍ�8s�du�`�i�%��<㒷�ř!^:Kד��\�p��~�O�|�2�rԠ��d����o���L� �}R`M��M��G^�ơr���.��7�(�B.�#H	C3(,��z`��v�vN��X�*����m�2j��G3����^�}��-��,{�Lw�_q P��8-�cߗ���P�>�A¨zg=�z��RKg>^�%�͖*��Զ�=��]�����嬇�/�}�8N���/7�Sm����*�^�+�t-_&�ů6��J�U�Y}��]����+|�*���6NU/}�λ~�F���5��~�EpԴ�\񚡱�ɴe�A�C���m$#�ݼBf�ƃAb�������|ؖ�,:�TPYQ�J��bQB�oN:_���"Sym��ܝ4���2���KM�H��N���~�[\~���+�dO+�r���rM�OU(eΙ�3+�bR�voNi���R�ks�|+��A
��7�1C+w|'`�����aɬ�P��H�Q!��;G)-�%2��X]�jʰ^&��m��{�V}�~��d�+���� ��d96u�l�|hi=�i{��Z��~���y����ޕ]o���Dԅb�>���z{'�B�Uo|������Ww\���0�)�F��p�l�@��X�C�Մ�ץ�R3���2n=a���<�+:�:�Sm�9�����]]�B�{��g:��j	���{x�p/L�vsL��o	�w(�]�>bn9w�#֪ה:��0͞�����0͓�\���%[G9��d)������덶���=�4��u�9�쿝�G2/)�v&�2�t�DB��'�%���4l_�����T�˪�6���]aU1�Gb)c]���?�>��,)smB��Rw�>��_Kl��ŗ��ñ��-J�=&�u�u�/�Sf�.�],�*�p��y����>N�f�� �B��A i�4�^��d��r��߯p�x��@���S; w��;Y�.��c�3��R��4�([��'�m��U�0���\g"�2�qq�м�����Пp�]��z�䣚-4Ce�i�ER��4&���)���GCY+3:7 �]k~��Q������o��jO��~$׿�C�mT'��(�|;�:~��jf�
��>
�[�Ѡvu�.R ��#е3�4��}.�qKsU���>�Cᬃ�9_��?����*�4:7��~\�q��ԫo�>�C�V�C��6��E���S�U�f�k �5���u B��({�➀ӣ���`?���|F�h��
�`@�kѫ������&��5^�����p�G5¯�s�&���j�V �<��d G�=����%���ߪ�]��ZY{0��]����	��9\���U_^{�	�X�:Mc�\#aيrF� ��m�-
�,��h��x�Eə�"�	|�D����F(1��'��u�B$3�8��c5FE^���^��P����ԑ�VP���d����8~�3���Cב��NFT�C��&���VAf @Fi��e�0(��Iķ��ghe������=w���ȥ����	!H�خ��t者�8g(M��=��^���G��@�cS��j�Q���0��)�tD��ܲc汀�瞈�}EcS��nR�r�i�O�Ȅ�P-YJ@u;:����݄�!ˉM�`=|J�R�aP��~ێ��d��B37��w�A��[�4N�qVD({"}_�U���/�����:���I�	2����\��m����?��p���$t'����hȑ�H�5��v�U�K:�����@z&�7˒7N5H�Ư8*N��^�a����}�����\ճ�y5�(�a��IGnQ�[/�7]��$��k�+!Z�;W�&�����T�;�<�v��a��:ֹ�p�����۾B;���-�]���[��K:���m�T�;�_��e��ƿƒ��p5F�{����;�i�k�n��59�S��X��J�G�VD��ă^
� ��&t��9�g�f���򴯢w�b�4���w~���h�!zߞ��j�c��:�u���.��ei��g{��w��wn+�'cԉ����;�aA��^�OB��aT�!.\* g��{O<�C���J���L��c^=V�њ{��M�g��S���)��w���5� 7�eo`}/�}8��V�hTYٮ������g6��p��k|�:����$׸�<��[D{�(�aj��ѿ}I[3�p%Y���[h+�J�@Ն̮�.U�W���_�)�r1S/b}X]�7T�x-����-V �GS��Ɋ`{���;����B�n��l3�4��2vC&��+��50�鿣«�K2U�7sC�Y��>𢬢N� ''�s�c,<�,���1qJ`}M��_U���҅��=��t ��5>��tč��=JK��j�.jF�yT�:Q����X�6���Y��o �e�d���F���8�C%*?�0�� �;X� r"@����⬹�6����1>]A�vi��@���&a�D�k��X��p�W���1�·�L���=(�J�2�z���|Q���W
�z��M�\�IEX&�-�,����(�A���VM=���Q�10J�����i��2�υ��x��#�k!��s�=�ۗ8�yy#�j�܀ʅ�15m0�*[Y𪐓��L�3�"�Q��ΚES�Ck��i�����z7 ��dz\7K�q�5@eB�J�"+�1��l
��"U�����0������)�W���H�w�O���TF����܏v��A���=͒�y")��m���>\���^E��oX`��X��_�/D��h����3祦4*��=n�?=*l�W8[�RؔD(���%��b� &�"ApF��0ď�DB(}�d�qG��í����ہ-��g����n9���?��V<2*j��&rDŕ�>�pB�!YAN�)��0��x��?�`�e{ ]�*��d��q@��1o��A�>f���s׶ЛF9c8��V2w^�"]B^����v�ZO�ݏ����w�)�}b����(A_�r�� �g|8��x�^l���4�����X�0�|4��Nw�0�ms]�:��QH�	�N~�&�Q��[a��h�C(��p$��:�Ed�%}���VN�a�\KO����@�53iע�?=wDB�m�
7xl���(���_y�,8���b䔛�Tk��VG qY���Hyƙ`�V��H�e��{֏o��X�6�d����+��]�îN�h�a�==����Pg,��b�a���	5*ǻù�<�i�5KdZ1s�k?�w���@�?&�c�04�BzP�DH���	��������i3ǜc�mī�Q�4�5�Ʉ��h�Vo"f�q��YY�YPж	K�*��_�!t7�Fg�v�/�M3$���^HΙM��U�5�Y�e���ń��X"ʯ��7,}Ø��Wjt��$�ݕrۅ�itapr��/F G��+���R��2tW�xZ�g{]9��Mvz�PX4�}H��aJ_0m�ژ�zg����		��gR
|с�����c
��K߹�d�>6����6y�y���>M�=�ܼ��2�jZ��r^�3�x��O/���X�.j�U�³n�$ø�rp+"��4KZ��ĺ��\�ʽմة��n�U�����l�T�+W�,:�Y6����/�Z5�f�~�/�8x#�,�/S������?��b�����mx>�j2�!��Ǖ!��_h��=d�is{;9�-����I�ɃM�Z��p���J���0��F���G��>�-�5UO{�r헙���֩Vp�&]�?�"���QМ���ѿ��Q˶h��e8�gE��)��	y~ɠH^|vo��Ema�]�hw�7Mg�M%�S4m�w>�b��#W���������!1]=)��$���E�s�Ꝑ�E��22)˥�$�	Ox�o�O�~Pd>�b�z��YH�I����Ê&��S�q2��������!�����GS���<4��K������|��Rݫؤ(�\����/,;���Un�����W�H�Ԝ��c��DU�z�|!~�+(�9$x
�׀Cv��-�Hp"��`ϓ&�F�a�>�<� sHw�F��Zfztc��c/�v.��2���ק&��Z�/���&jޜ�_��>g�CJxmF`�`�c��z��&�	��ݔ�� f �<ڛ��Â�L��39q�psۜ�i�Q >��LG�W#7T�A�@��#�yH�� ����N��2�&�Q�����LB������Stu��{K�����*�D�̦��B�%sJ�͏v ��ܳuuex/��e�gxoVrҔ�W���o���h�m��}� �2/c�^8d�0�6�!3u&���z���ް2T^���>9J�J�Mo��B˃�@}h�P
�N昪
��M-A�3�V*e=dM���		y��5�b��PE17L����J�:tFZQW�U�r����
Λ�Y�'����4'Y�T
o�5�b�����D�nBD:2�<Bt']󀵔�-�uCM5�]�v��^�;�yf��R^���E�$'��^�z}���-��cI�m�\�y��J��M|\�0h%��(2~�b!���M�. JT+�FJ*���$b�������~����=)���䮤�=�����?�\4#|�e�L�3������[+�Ŕ�W!�՝y_�L+B^��:ɉ{f=j�{f�֔�f_G	<����/[�O��{�����ev׮�:#�I��IP�wk����%%�$��|e����y�F��d	 �ȃ��Ҷu�C��!����?��*�`�h-6�*v���.-يK�)�� I�{q�K 9�S8�w�����ѿ�!�C�@q���&�0 �D�2�iװ=ո��Q�:&D��j_��;7�E_
��E��_�D�4O|G��1����_\m�A�\�ܾ�a��S��z�W(�7䈐�Ǚ��AG121�4��끖#'�Ŏ7�Oad�$��-���K�a �'���\� �&��V=Y����W�٦R�&&�|��z�m |���)�T���;�Z��X����_jF���8|��M�4~��:�"�
�����Y+Czu�ئ��WR�R��X4�ƽ��;ַ��X� ��{��1�\�Qu�c`z��EN���	^q}���kI>gZ����_�tIW:�4^&+�N5�^K���Bw+N�׀����}r�~ ����A�VH��#��z�+{��T ���D���'j�-�bu��7#�@�Sz�+
�Sl@țb$d�{ˢK���=���_�����F{HFQ]�i���QcE�O�����	}�n��qC} �,q�\�\��*�#�� �M9�3'	uw�ѯ{���3`~|��)x��:�u��A�p���jW�^�D^߻���+�B��4�m�dJn��>�/X߶F�7w)�C�8!���J��VV�5�&��m�������������8Z�;M������oML��X���k'jv�~vQ�̘��d�|偢'"ʲˏUz%Qht�_�>�S�Zv��}���`����=`�T���L6����Hօr}&(h�ד�G����N�ѳc��*��,��h����Mq�����\P�+��3:ws�c�d� ��;�+`�O��އ'֚ͽ3�A��dSU����;=����.O��3<�R�����R'�2��_/�|��z�_�q�<�1�S�$�fZ-���蓤�����ۨUSڧ-�q��q8Gߑ�J��]�}QO����$���<���G�ܡ���q��'�o�Y'	�~�1~�)v�W!�h8���yr�[&�w((-�P��Q����� Z?��\f|��GMs�ߋcB�|��-O4���a>����*��9(�P.�a�m�����]B�ͪ��q�,�Q���ۊ
��"&�6��G��M�tB�J�h0��E��Vތ��"�A��v��g_�h4Np�B_�6�D.-C��p�v�i] ���AX֒�]U�C��	��N�4`tj�E��!�#����@�4��#/�L�~P���:��٢F��	ǆ5�\uu9�zĿyD���d� c���&U{FW&1S��\��7Pk�/Vjģy+s��R��Y���8�)g�CW.vmV�3+�S�!dC��MB��N�-�=^^%)�ί�ʈV�63�4,�p�P�����z�����XY�H[�e߿m"��F�~2��	���z�;�1Z��ڥ�u ��w��A���Q�,�Z�9����kђr���c~u�u�x�3��bDUv�|���qi��q���$vї�������Sk�7�y��<0*Ds�}�QO!��
�̰}���n�ZT�_gL�L㇛�I����qMݥMX���k f���\鳎�K��Q�τ����d���^�hΰ}{œ+�`��+6� X_
YX��k��
�`�V�חH��

a_��.��x5�8��'�s;������`x������W~��&�t��5g���E��\F#^U���P�c����Ւ4_�	Hi�>H�]Q��G���]yB�g3�-�V��"�-�?Tę��X�q;?����z�����{	y�$�rVܙ�M��R@����k����tzȎ�t��&;_��@�%���=L� ����n��nS�&�Y�(K��UF�.=�$�h�$���~R�%��}|@{|�����/�x�*�g<�k֗�{LAT�#��RߣI&3��ț���#���k�l�>h����C^4z?���1:uD��Q����N���\�����Æ�?;���)���W�&׮�V<5#k;�)F�!��$ny4�@0m�*w3S��F�tK��}�� R=.x���~M�I,�g��ѭM�&��:�9�>AQcZ8��� �c�	��7�j�� #4+[�m�p��pfȂJ�F=ʀ�V� �~[C���a��3a:~Vb@��YJ�0�6�e�i��0��t�Č.d�HwaT�e	r�v^�'�����H[�l�2 ��Wa9���2q>ۂFW��!��K�)x%m��������EN����o��� gE^ƊF�D_�
QaHF��!�E�4=fa������x����P��|Z� ���N{x ��1s���*;�Ga�,�I��u���nȪȺA�b��ྂʧ~���p*�,�Ǵ*�_�-1�s�t��`y��H'�"FW� ��Ĭ�v��<��ߕ��zzn7�O��ֿn+v�v7�z0�T�Ec�WjU�y+l5���je>v`�'"oiU�� f\��1,�R�Նd��W���6Ҙ��~b�<x.�4ݞ�ʶ�| y��� ׹*Z馉���N�������%B6 	)W�������V�+S�1떇׻���nc4XK��t#	 ;�oHԝUAS�ݾ�f�/�?�����?f�yg�H�-�gt�5k!��7ٜ���j��r�`H?���G�o���G�'�}�U	�e�[�O�ۦe�(�$WZ��x�H�g�N ݆�1w�K��w~���PY����9��eY���d�c�FBȞIh����'��# ���j�BHQu�6x�&@���<�6υi�R/��:0��羭'�hL�O��n�����R�0&�ex��6b�VM��Y����*����ފ'�$������y��{ چv�G�k�șj�P��l/vil�/>J'V˟S��5��o�����ݔ��QUE�)sӰ��͡���1a�E��E@��9@��M�O�K{TъҪ�-��B�t�z��n�G�jԫR����\ɗ/#�6D�I��xC��4� Lh�A��	������V�fN�@����VG����@���%vߝ��Y�K���?&#gh�^	yN����I>&Hb-��[޹<�8L�W�a O�tk�,X��)~PL��c�WI0ﲱ�s�6�hMz8��R�MQ���յMe
����<�>������u�0]\��x��'���@)�h>J#�Q�PJP�֙M/����!��Ƒ��r��������4F�Q��K8��c��l��X��#DM���=�V6o}uQa-��q�p�����X���:�H},�Ȗ��܈�u���rG��Ga�!�3=7o|�����0�׻�\uح7<,l*���p���e����/K7�Ƥ�����H�NrE)��������K�A���s��0�t��XD�oy�������FX�O�t��)��Qfcti��W�P^<�"a�efRд.Z���X������Ǚ��$>���&sZ�����$I�AR�Q����
�b���e�.z�]�!?g��	}�(�{�Vc5��>�D@��>��ZϽ��e��~}����.=�t��-���Y7m»����]�r���>t�Ӂ6h��!��R��������Lo�ޯn�D�3��t��l��B�s*�J��
����ѥڲ��L���-�/ �AKA��˜\+QV4��.O��qN(c�J�T�P�-ek�<hK)w|��{�5�ȈL�z��B�KK�V��5��h\N�W��6�j�U{�FNE�K�W��J�3��a7���Wc�=�I�Hd�M��� Ӭ[�H�YP����X`�Fx�Q�2

Fa�id�[�]������hJ	l����Vuڼ4ФHU�I:7!�\�!���t��̐'�m������7f���z��2�(��-��W�wv�|����1�HCe,SeG���\%�#���R�ܠ-��M����,�[�yT!y�v�[�Gؐ�1�3�f��5�c�Vۿ���Тa��#��
����ߎ�F���*a��.�j.GK��D��.j��}��|���ŵ�a:������0o��E ����*��U�8�=�����E��dM��H���x�8�à*��h+O[	�� �K�x8=���0|6c�l�٫�s�U*�F��h>.��*��'iW[t��rU�~���;��*&*���@���2���.����9x�)�~q�A6��X��';�%<(��2�y_�R1?nכ�I�՜ʻ�L(��d!�� %������о�S���8�#'V̾(���7+�=��?��)��"���&E�$�>D��� �Z����:;U��;\\%h�s�@�/k��4��dz�ܼ�7\���.VE��N����������h߶G�����@aǉ`�E*?$F(@��oZNt�����)�D��T�5�>:��[����vY�ޟc������|�!�ibht1��2��C�W�0�h��%��0+�j���r�9�n��!�Y�/��d�do�-}����������Kǽ�dc��>��0>�S<�ź9��9�������]�@�%c��>��< ���v�34�l�@͒�+���.�22s���Ln��+��1������+��l�w}�?����[�E���_�����z���%��'�U�TX9�۩�g'2��Ò�T7�,����+�����_�s�WW�TxI�0�����hR] ,خjʄ�6J������a�61+Ҋ�D"��5B��R׋�uf8f�6$,]�ݴId�gpl��5�(a�q��d��N���I��睕i�#f�1*������=C:Ij���'���ϛ�gDʥ��l��|��JW����ݺ�xȁ�SU]B��M'�kګ+�����
?�raѢ ��祖p��dH'39 �]���zg���ƥȳ�s}��%�0��_�
���i[H� 1��Η������G�SE�gY�ܥ������z!kC06c��Y�J*�B�=��o]�����ϳO��2j�W\����*>�q2m,�<���0ƙ����jpEF�����hK��)�_oV�]�l�}�՜E���H���mj?���v�R4JR�(�"h*Ag]�߲�����G½���p�b
Sӱ�NltC���j����T�/}
��;�FDR�3F.���}j��p.��?kr��	8S�\!J����7�$�a/ڳsc�j��*d���@�[-j?��:n��]S�:�TJh�``�F�l�V�0�����4��BVW�A� T~�A���4��՘v�)�D��7������l3d�����Xn=_~�Sڵ9Ʃ��B0O�s��\7�Gs��ʠVd����L_K�;HRZ���J�7�Qr�R���g0��e�/pں<�N�D��2ddw-Bl��� <���}`�ީW&�bx`}\ji�\2�'�6Sk��'���G<�����H��y��T��ZM�Ӟ�h ����F�oi��C-ԛ����r+?Q���YsKV�CO�vX3�$+;�9/�}�_Zض�t8j._��s���⻻<+W����"���?���#_Y&jQ,�~izŤ4��g.�%ָ�q�hC_�\:ײ���aľ�\��ݨ&�<c�R*��%�g�=Gt�B�[ ������/z����S��._Y;��O����Y�IGkhp	��f�8@���#�f;�w�ͦ�.�'�ȡ#p�ep��SN�jQ�C56.�A$�l�#c�[����v�4)� ��T�)�����]�'���lMRU�$�R�=����YO����.�X�RD<���R���0<��;&]�"Bh�}{��n��1��<�`�^P��lܾg��N�+��G��8aM@����'FVX��i���۵������R=��'���Ȩ�Z�����Q�װ�0xr�a	N���:��z�d%4Q+�[�s�$�V��LI��	Γ�bD�u�Z��a�������V�~T�#/J�`��I/��a�H�0��%J���!�{�۵�x��_4 Y�̃�ZB�H�:�*s���QNt�����f��?rV�P����j�g�,, N���������j�(�W�I��E����Y;�%�iq�<�M��*yaB_Qe�XY�����Iy*0�Z��[dWtD�����b���������~��V�E4����P��ϣo�ڮ�׈���'֝L��}�e*�:��3��ՠ�.�>Z���>! �v	_�0�6ϴ��#���D��4m��Ś���/��)q�w��#�є���M7��)�]CK{�M��aVQ㥳Q�5l&�+�G]4&���vf�ȇ)`�� �;	E]ƍ*����e��H�.=��x���c�a��=���ZU��>!;Hm�XR7����x�~��k����G�&���E��e�����R1j�늢�;�I@4e]MU< ���!d�o]� lE�aޗȗz��EF#CgkR��?�cC�B�\00螂��o6l�O��Zk��&��ZGBIi�f#ʄ��䤎��h�Gw=kD1�,�P��8�5;'��m����,��M�U����0�WJJo=fc��*j!D�mh�׉��m�lWz���e*�W1�\S�]�o�Z�f�Ў�̓A#�
3�v�lN�_ hb�;��%h�K�+��;\4���b��4ʾ��zK�Mw*1WT�:���}�*H��k�0IE>��p��$��Y��7"���M�Y��������4�nY<L�Y@�Րh�BV�=�N�hN 0L�VqJ[sj�2�(R�6$<�i��d(�F�'�3�R�ݾ��Q�[ld�� �Y˃h���8d������/�_�$�_!���5x��N�~�W-����b��P���]ׅ��f�$x�y)Ǥ<�{ � ��8p<�V��?E�c���K�"F�o��1'vE�wE+�����eRɹ���^J��W�~�<�\#7p��W;����D䡈L1-�b��h|7����y�Ϡ��(�9�E�bo��`ىw��"b��{SS��Y��:��İ��WP�}rQ_���K4�^�C�i�Z���BKs�
���~ј`���^5�}ʔFf�b� ����V/� X��E����԰����]4PW���ެ/y5���7��nH� ��ėm�Q���