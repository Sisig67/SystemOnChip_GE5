��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���!<So���2��E�!�7���feI�R�34�F�\1uR�XO.P㤳��"����(W�����Y�us�'�V6g{���/�Y�^( ���Ne�[�����8�1��{SZ�k�eZɇ�FUHn�i!��Z�CZ���X�n��U�tr�Љ��������z]O������փ�=X�MG5�G����C��{����a�}�C�Z��b���>$�����z�[��l�;o ���'�����.���%�1k16oҦĘ>:���Ai2�L��������
n{Yt�n!������j�8`��Z>򴒈t�RJ�^FWwl�*�GR,�a[��>� q"��?SA�u��	P��A�t��A����}�R��Ѱ��ÿG�<�=fH��;��?(��ڞ���ăi6�-Yd�4�>���t��I�[օL؞�ܛ�ZN��<�����J�ds��#a�D؏f3�/ݕjEp3�ļ. (=�T�|� ��t��O���	Fo��8�05����a�{�,�-o]m�|q^�ᓉe�5H6��4�iU'��?��>�c��G�B���+���)�p�\��>�1��Yf�kn�0B��UR6�J.���{�I}*}��B6�X�tmi3 ��^�3�	��ݜ�T�e�h%�ʹ�&�#'�!E�!U9�<��o���q����W���T5�
%(�8���>#���~y��8�����t������iG�oI԰A�(���|6��vw�t�'����Z�р��IZq�Z�r�x&�|���L��A��Q��0���:��l�`���Z8<X^�I=~����F0
R��pȄ�֫p�|�I��B��6k���sI˱��)�6L�A�t��G �[l�8"6_%��NY�v	̚+Kh��7� ��%�+�(+������|�%r�������mO��Rշ;����>6��#��t����� �4)p]�3��� �Tʉ��5@��E�������ǃR�r��ё88���w�I$��h�NU w�'�*�G���h?�3�>΅�_�]�mr	�5��¯s�aA���w	��;��g��7��]kÚ��L�^���*�~�Y�艂�=宇�5�]Z��z苪')h(�9�OD���lUdP���PPJ��I�	!�1��8�q�W��mK[��U��h�|
�WB�T+X��mY38F��0����/.�"٣�^&d�L��P?"G�F.<�����1\Wo�/��R>�i ����{�=��M'NЎ��qW^v�7��sՖ#����Vk�..�	<oFz$�g]����	�*�(m�C �G{UW�R���׃��Q�q�^njğ3@�>KUuT�n˟���=K�Ds��tߞ�8��#�̘K��oe_U�j�T�l�ί��$zP|��wJ��c7��_I	[�~V�s�Z���g#�[� �� ��L�A.i�.�����+�w��z�@�A1~�x�Q�`��t��Hh���#�;z֠R-�����K����>�	J9�q�������QC�=��3�k�[EJ�;��\ӫ�?l��c�s\�j�$�)��xu�8��61,��v�F���o�92��`�H?��e[DOL�cF�]f`�R��K�B�ԇҩ<g�&��{=��a�Ƀߓ�;�)��gp;�R�j��.8b�L5z��E�"���[t)�瀱:��\�󈑫�|�o2�|kF��Հ��l1Q̏���&Β��K��YD޴0ĢF�����S�r=I�9'-a���һD8��	U�D�䥍5����2 IT����?l�6A'Kx����~����	q�m�}����!��sY0��dRK�R��?zZ�K�(����c�+U���j�5�����l{%c��F%�;��xTڿ�q��N`c5B��"?���1��r:�԰�a���h$/绱vi;ZV�mb�~�-�!��,X���%�n��H��eI�����	C�o�Ԁ�i�9?��1�lp��裺��L㱳g��귔�IA����aX8:P6�i���9��
�oV�ig�uP�,�
��Qݞ��YH�z�[��c���9.j!�h��y'N`̃��Ӵ��Y'�#g����&P�����jb�5l}�d�����5�姸c�,�l9й������Q6@z��O@0�U�2R��o���4�i�;��ub�	x�k���j����E(�|x�=r]��e���^���ph�ܢ���*|M���6� ��������n�R����|�׫H�4��WnK�����3�ಜ�
��wET%�|A�|'o�8���4�5)o7�J�'N��'��@h�`Ԗl_��0і�s�UP.�P�!~B�����e��躴1�x��G��dc}|�x���c��H���tq��iA\#���uyB�U��9�ǆQ}�q��e��h<O:e��������������=T�(y}g���x`�C�!��8�N�DU {�"C�e=�Z���L�ʅ��j�i}��F+:]��d�D;��Nq�R"��S�<*��gu` e�{v�8$��_SAnR����dZ�#ɜ��q����7��ӗ�I���W&L�1�1�Եx����3͞hhYXnmKŶ�k""�Y��j̒�z��@^E�ۙ�n<�hُ]/�jo�+'As��o"�+��9��^��kq��:ͨ!jm������#��'fF��|�x���@�$�(b䤛SH��A�`]#���$��r�}��|I�8~���ȇ,Y�O�	��1l�X��V���ufB�^Mm�-cJ�%S T��a���0F>*��N�f���d��k���pǯ��-��JY�HU�E5�$r'��2�QPd�`�<�Lbݶٖ�x(��M�-��ؕk�#�G�z��BD����n/޾����z� -�? �v�`�~���h���[�V˾��Gq� W�y����U�DK�ɵ�ܗ=��0�K������enP?
��2b7����j�e���:�
�&ʹ��u݋��d0�	�)XH�߲#��q����M�{�� gߏi�M���ޚo0����z���Ϊc�L�"���V�v�����{�O�Z��O��ɚ1Q��F	x�� ��
�.�H�}��sN����y��;yu-n7�xe��,���ўh��f�o_"n�j�OM31�Xi?k�Y��0�nb9�B$j�s0pk��%}����=n�Ĺ�Y�9�^T�\�1 ��V���N��_������3�U�����=y����}��0@/��{)M!}�۱�����u���Ǆ�c��p�e�M��?#�>�U��>�t�cSo^��^�g���Lh�Jm�)�4-�{(j⺣o���=K��O��!�Z5:������7�7�����ζ���ЋǢ��M�|p1�m�{8�d~FU�d���~t�j�^�d�SԷJé!�����57�b��h�iJ�X�$�NoeQ�r��	�?���KFl�ܟi]S����n�[�'p�NZ.�s�.��������_��Fnٍ��s���eѶ�&{n r�QL�,K#B�pr�������s�jр#j6CkW�DgGc���jk��5fP��߽�2��kW�Nx���>S.'9�������D�a\q�y;����R��ӣ�I��q���jr
,S}��������H2W�e��l%��p� Lg�Yԧ93�?-��MN���9�>��˜p�b�\d%�HѦ�8��ɟ�w�ub5��p�j4y�����%�"уL	���
 �D�%�����]�)�y�$S4��F�5��u4lW@C����p��M��$��B��Id���-'����B�㓔��f�� %������z�;�"h�fJ�^u,I���h��'\��ih�0��Aּ�	����v�Å�U���.��1i;��A�����qܘ4>�[��?1"�%�|��]U$eI�f�dhD�^p��l�yH��^ƣ���#>T��ս`	�>�ӇW����c70	�dO�C�<�+@��{�����*,؏���յߙoK�sCȴY��K}����4���(�O�	^�NX+��%ߵV����.�w��5��_kѩ��k��UM�B��)LǮRJI��P���+#�V�O�-��/�͘�ykߜ�gm�%ۨ���w!&�s��Y�WHo�� z�x�_W'T���%8_	�,�]2���	~�֕?nм���e��+5؏�%���d*��1bOQ���QN/��"�/	m��Lw���i��vE�(ro��������4DxF���JE�u�)��t�{����YG!~���s�A%u�,*V�Sp���;^l�|p?o�ԃ�%J���͘��ܛ?�UIذ<V�h��j��R٫F��zJ;j#��j�����=F
��b�`@�3�[�[Иa0�����mnL�p��7>�4�fB4S�>����oD&p����W�b�X����}�s�7GP,1�n�w;��ڔ:Ջ��I��ۓ�{�U@؈�͜�oT�V�jΕu��U��ʶ��h��<>����'�=�h=8-jUl�����k�7���!�6��y�ɺx/�ᨉt%t�30$�C�\2�]>���7�P�E��#��i"�����%{L�uה�\���p�b����`os|�!�M"�"@���Y��g:��NZ��$����k\u����~���VO���tݞ�����x�05DI���G��f�[[ϕ,7��ͬ}��YM�mc��2J�� �'��-kQ`���l�HYo����=�,.��1�h|��>���4��D���y�'a��z�Ks��\K|m�^?�߮	h<��Ӛ:R׀�n��O���3Po{����K�O@/�]�ϑ0#��f��kσ��
 �/�Z+A�X���n�!����d�_�}�22z�܆��ѵr�&2�9ҟ�����#_d�lg��ڮ?������o�aT(��m]�ᵬ�*9�N~g��]����>j���h���T�����o�q�Xcę]�������ob1�L�� ����E���g�7��Tah#��ߘ�CN�����%
/����Q����D��bC�L�`�4�d��I_/B�~}��9�!7�ϓ�y��������3�d��Gj��^e�38c|�J�Y_��k�F����א��cHD2�kY�|Y�-!;Ne���E�
�{-����G��K9-&P�vYHH��?�鋊���P��E�e�
>�gA�I���v�[�=n�>�8=�"��M��"ڤ�tޒ�Ӹ/r�HR?�T�`��T����?�ۘi�`�J81��0Q��;������ف������ӊ#���>\���$J׸��'�+�-ϕ��)_�C̜�i��/��??��VKy7�y�w��=*�����Z��s��;���w9/EGY��;��K�p.U��� �L�ȸϘkA�,��ͩ��eǂ�L��;2V��B 2�H
a�@C�P&��.�z��`Rwƺ-�I�� ���2�8�X���%1;���P�5|�8���א���E���ǐV"=J�2��/V�3<�C���N��[X`CG꯲�	5���M�"U�.Jc�G��U��5HXzL��n�����V��	E�������ipO�dJ�I����P'�tȜI�w"��q�1�y����.�X}��Kܟ":�Ov����x6���b(?1,o`�T��P��J������.197���ݮ����@J����3f6�r�=��;��f"e��`��J@��M�[ᯢ��3޴Lm����I���Ԗ�G��r�l��Uڎ)�Y�}�:V{(�ʨ��T�h��?]�B���j�x�Dy�p:�Zc�\sǆi�Ӻu-��<6C�}l:O�i�T��������)�wݧ$+�#u�:��P?ϗ���q��μ�,���i�9������
;J(�G�XB����*Gk��;(���P��IO=;3D.��&a��{Di$������B�vg�)(�ᢧ�N
�o�:�$�{��7'�_�����
3kEf�[���g��D���M�A��ƕ�g�7��#�9Z
�+��m����mt�pw���M'��\|��z�Ӆߍ�mP6?�G+�c2�m[�4���N���F ���pKiAᙕ�g�s�p�a:ܮZ�M߉k��Kϻ�n�r}?]�F�a���+]�9�5W�b;8X���SJjz�{?J
��t�yZ	�ӭ�2�<K��;���L$
&��%q��'0(9�877M	��3sG������NU�U9 *��h��T+!襈)�Մ\m��a>zd��4R���ꛒ�I��b�/�D�B��yxo�_��1b}�,8.�B:ꪲ�M�F�����n�E_�M^]lC%�1=�,�f{q0�	unKZoM�6� �9_n�~�sTZ�/=8
]�6�q�����ǰ;���+�,.8��*��p���Y�����6y��(ӷVB"^D����WX< .pi� �=S�k5м�9���.�jK�rJ��^d�	?
=U��5�R���_�B<^N��4�L ����F��tB�Y'�D�XV�vF��AQ���Z��0���0��	��rf�;z��B�-��_.Ĩ߂���W��[��b\�G���w�8�$��<��L6�"��f|s���vf��k[�m(��|�ú=�Ǫ��9�!vt����h��b��Dc(�2�]6�\S���ӳD�4ξ߿��I���
O=T(⥤���k�
���"{�7b9�z���*�N�n�)�	���hMwQ5%0�I�Yp��nQ� �@�������p�Ar��k�H�sp��y�)Y#�6�a�~�E(�@�dq��[<�]�y�B��5�b�{{.��嵶T�^��}+S*�PhBL�&�%��]F'�^���l�w�dE�b�WRD�
J�rC$y�<�he�'�d|�e)�j!��O�h�ǋ����+Yv��.s��p����p��u�/���C�w����ȳ}�w;����Xr�����l�Z�N��QW�Я��E���u�^;�̻�F��4��U�%Q���GA�	;ȑ�ڶp�9��E�[��U�
+\�R�чf�����r��lCk�n��l[H�o�D���+:���j���3|�`gJ=쩫C�7��Q�\홞�(�U�<�q
`d*΋��Sa�B�q���nPV�>oTl��S�FT�=�ʫ`ť����3Տ�	��x���3=�����}��~7,u�u���G�E�iJDq���p�o��~�NK���`޶8%�w*�f3:�t����nF*�XR�`ۦk�=1��x�ôd��������he�~�kkv�=4��ҹ@Jz@��j3[%۫�П?�()�U),�p�<�I<݁�_><?��F'��a�O�EҲ_Uҕ����9wߪ�"D���ӹ��Y;g��J'+�]'�c�S�!�S��u4�j�v����wSLv���o��l�EODe�(�E�ؓ��	�. �e����i��I��b�Ӈ�YV�-;Q*˛]�f<��g��
��z�NQ���1���a$���ʇ��A���Y��'��kd��rY����&!��!�[P�����E�{Z��M)��X�R� �9ۂ]����p������_޴��8'���jfk��9IM��\(�� *�׶�c�P/��X���9���B��`���P±F�{�M�M���-M�����!5�G�4�����զV1�u��c��j�zJ�	6#V�n�gd�!_r@FTA͇���w;�?5�Ɯ���N[2,��
TH�fk=�,{���@;���B���nɍ�mV�tը�p32*	�>�b�t&�7w�iϙ�x��-�]��%���D�mЕ����Q<n���� �\���O���d��3Dh-04��9⟁�>���M�������:�!{��5���������}��m����j�4۪74����/'�o}W"DI�=��mW�Q�蔧��'�b簳E�=Z�P�$���,)H1����K���x��s�W��k�QZz��)���䋙���J?�';��+��)������0p&$�� M�͉�A_3a��/\����"�B<N�&��0\�L��I14�R�8&�Zm��4G����K�P[i�a��u
eY
g�B�t��i�� �)g��ͳ�o��}���M�S��l���@9j���*�<�#V�t��y5_�H�/�G��'f�Ҵ���[��7��rx''b�%r�����<{�.��)7B����@m��������8�&�ً
�y���ė�R�ɡ��|(��-�|���R��!��9�}�S�����C�傼���K�+�T��׮]���Ɇ���RI)�(:��@V�}u�5pt���]o�[�W�<�����B��#��(�Zq�H��^���i:�]���^��i� �tm�s�<��},�g��}��Y$$�$~��a����w8�@� �r`��m�(�0Kl��*��? ���"�}��w�hj�lU�����
D/�K7��L_�ev�#����hw1�J��W�u�����_��h�"[^��.��Hf�$~�ksj�Q�+׽���8�A��S��}^���GF�B
N?�ű��O�S���P/�*,N#�Lx�����7�H���4�y�!
9�_��#���!&lt�|V�}��@Z�q�E�rf�D�z��i+*Ǥ�?�cV䯆�6o99`�:�/HG���ӧ�f���_A�� ���@	��~%?��Ɨs5/uIhhH����B��$7'h]풷=�r�v��(ZsP���Ӥ��hg��˪*]�b'W�BV�?�ô3F�!�5�*����r����b�x�K97{�`嗲v$.j�j�ox�(�f�D��{Mӹޙ5'.JgC/�a�'�3]s���8����{Q)�x�mT�L/���3=�"�m���s�"Ȱ0�9΢7�}-�e@��g^�I�D7�������|�K�ì���cE�L��-
%G���h%��q����4Y;��p��Z:�:�3q���x7A�W��>g�e��Q�v��x�]'tɲy�T{�lAE�0�%��ӑ��rW���I|.�TZ���m��Q[ӻv�RO0�:�2u?5S��Xۆ���ti�q.�c�r��	�+��0)X�^z�󔭃���>G�+-�/g���g붓�۱�M��JP %��Y4P�m��(S�7[�2�q�i��_���o�׿)�G㾁�����|�w%��(��>�r�h�to^�Rj�k�&k�!_�%ՏM���oR��$��F��#X��G1���*��.9����.Y��)	�;�u�Ajz�#u9��n#4� � ���++F3���RB���J ��}k�g�Kt�b���xr(�$�V�)}�1�X�[�c䒮l������ְG������\�G]�x��4��Y<+���ybv�ױ̪��\�X4Q� �����^���Nq۳�띲�ՊT�~F���l��3J���r����C�w� ��Y n�B$8��Q�犌�'d"�y��B�v��0C�������/�n����h��T��h[���b ���>�$�]	��<�9��O��)1��%��4C����a�	M��Xs��*N���l�-lM�@�_�N��jzä�&\R�T�'�!��ɶ�_3��>�� ��4�m�6�J���$9բ <h���r�Euv��v�}��������U�LtT��w2v�I����I��9瘾кiܿ���]¸������9����q����U�wHRh�:4�>7xe:�Q�����3�k����惠�����<z(�FY<G�|!�J�	E_���91 ..��ȀuVl��[�s�pǽ���;1L�޵U,�&�b�K^⬟�[��5�iLh��Y�*3b_��q.O��t'�5r���ORF#i.���:�`�a�/fkx]��۪�݋hNr�&�.�X�1<Z��b���Q^�f�@{�P��������'�1�N�����֬$tZ�Il(�;ЈJ�� Ax���K�����d}�5@w9{�8Vh��8��{)7g��/���e=�5�%�V�ZA���������޿��꒷ܘ�Ԁ >�#�+���?*�Q����XX�-�xNN5?,r����ܧpAn�$Kk6�N�P'�5����)��*��YOQG�lG�wԵ�e��g��,aV��X~#w��tXW�`��r�N�P��[�����do����#�O�\�}�/�!��h��O!D�^C C�����6Jnr�/����D�ǅ�P���X�{y>)/!z� r� ��(w)F��>��25��)��3�A�����h/�s��on1�YN���/��[pL4�]���>�l�VVm=G�yz�V����o#ƀ�>=5�&|mHw`m���ot�(�	Ȑ�SE%:me��Ny2��K{�H-��<�(�Q�� �r����w�/S���/�^,�V»5�~ʢ�s>����Yqa\����_�q�T�Dt�=�!�|t�[�ݡ��^3�.�U�*�P`���z	(,CB�"��n�9	���y׽�}�ӄ�����46ڐ1:�����,�3xҺ��o�YG�	�n:
�'±?����Z�&�m#�i��
�r��/=�ld� '�q	�$�� N..坯!z�x�N�ߟC�,��]��-����!��Xlw��ʁ���|Q�KL��v�����kgU$�G7gf���yv��B�!���T��jY�Tg�֋�� ����_ ����2%��#�^%�Lw��ݠ{ �w�j��0���)$:0�缌t���|��w����-_%��Є��͆D,oB1�eq��%�~�i��<TD�?�7y9��a�Z��1[/�@����ؘ��d4�g C�>�'��B~�.��0q�=���;�졌ZN��G�\'<G���ݮ�Qm.��;_��E
W�qܛ؈袋��ӱd.���(�H��6֘s��מ���dn�ē��t�����4$�����r�ő� �YD��5򮝟�'i�kDwR ����7r3�C�����1�@k��4T!3厲Z"���y��y�c�qE->-^9pTU,äW��|V�s���in�:_ö?���?���ȳ��Ap����4�f�����ϼsZWC�~��n]x/���zu|�yx?��|$~�bv�	�H��=��xrB��e*�1����ٕ�A�cj�OS����9�?�PL�Қ���T r�S6�=ƉƏT"�]@o��q���7�AܩX`�Ӿ���CD��<5��=�����,���
���n�b�v��c�u�+��w��п������E��B��m���r�
/Ť��*���J�8����'�~M�c�����P�<��wg?��	k��/&ANBy/��[Cd�/�kI��Ԉ��4:>��vN��7�5��cr��+M�"a`��c�F�$>����_]�����U>�X� �sNU�N�us|C>�֡MOB�����`?�g��S:�tf��m"aЫ�������л�u�2f��Зv�^'\�pn��Xb���V-����������ɚ�Bp�0V�	#��s:d
���B;W]{������k�Y�-�2�t?~`q�ZC���9m��=��G{@��(�d�$������JV�v�!Rכ�t�N�ް�*\���i.�����x �̍E�9Q��������<�������]А�P�� ��������p��D�߯	R��?��a�S�� y�U���O'J�#��AxB���D�K�܇�����j@&"]�T�<���9L�*�:I�Y�:[���1�'�n�r��f��v[��	�p��ÆP�G�4�U8���o�x(dh���Z�|��J�@�
�/�u��-�%�fJ#�#e֓�����0�E�"t�����2�y��9�ߟ������[1�
|X�he��5(�b��o��w��C�����#K���zF��2Am������{�0z�B��R?��ES�f�ȹ�a��W�������I3f���W<��1�?�ai 0���O�*pP&�����"�q���fͺ��nf�)�š!�V�Yޭ��(�Ҩ��|uBT�)�Ъ���ό��r�{D��P�"Fy��0{���b������ӯ��S�y��
j�n�6+�!�����1���$�e��8��Z�x���k��P3_^(�׉i��uW{�.��z=BaSdA��]%��?� ��?3��9՚e\��Ʌλ/"�nr �E��#��w(�[I	yR�-y��=h���\y��ȗ�gk� 3�"�@ܦ�=R
7�������']�Z�ئ7t��7�!/�k�#�W-���_�������ӭ�:�q�*^`(���V������P3"�O��b���ъ�f�yg��G��;h��8EY[bd�>m�A^<ĳ�]:��������j�V
������`:�-�I���p�+V����c���6��&�����ZV��`�&��줻V����f���ֈ�Zq�M���a��ߝbeJ�}@_���#����.����.q;)��[l���MA��nW��I��}���V36$ Q.�*]dl�	ʠ�������Ń�i��3!�g �����g���`m���8��ƒ���1�������\�J�+Ñ��|�9X�;اyKc�<��FN7�d�D�"�='��`�n�,�5*t_�mA+�s?%�2��������-I��_:Pj�+@|�]5���&Vy��H��쮠���z�3�m�|r�I��iP�i?���}�@cM�%hyp �i�H��lv��XC�DH���c�������6� �e�_7ir=L�w�����~��|XY�0��;Z��^�y��[I�~*{[�o��"�"�̻��h1߷瘤v���	>�Ơ���B���k�6��8�@5!1�6,]��=�T���8�s�}I,Q����@�_Y����%���aڹ.��c����i�@�DO����˧� ����
o��(����h֐fP�R�u5
Ҹ+�O�[�>7�v%�kNd��v�<�6���:��ûя�L�l��)d#��ڭ�7�e�c$�Pd��NS9�w��Z��byя�_=q���J5���l��Q3��JI:Ծp�>
�m����%/�
��h���S-lrw���Q=ef�4�a��
�ʢ����}�NȻ�M�v�0�Zؚ���$�p8�m0���EOnCIH��~�|�*���NR�H��<k��������0/�����H��A��7�6Bk'�v���#�Us`�ڙ�,p���E���4�.	����?@$��c��i�ʷ�
R�������Y�%��,*�5�εQh�~V�z�6����L�8�8LF�rSg����iǻ/|�K(�����G���VzʘЭC���8;��$����B���Q�Gn�.��j
*6�K�j���n��Ҧ�X���FI���X�[$tg��p��!�TO|�)�qf��\�md薪�e
Ăq�f������;g��ofJ����`}n#'�/�ێy�ై�(o�$?�	�h�`��I�a7�ҠEsNq�la�7��K��kɗ�]B�:Z�K8P@��ر�{V��W�$�f�L��:�T�!�-Y�X��,Nh��,t㌠34@X���@yC<6��r�H ��gYw)�H<�z�t���� ��x�f�q�#g٢Ĵ�"2~7V{��Z-��(�~b
>� �h���QT� 6ȳK��,�;P�� JÆ-��t�~s�
�k�J��CT�O\]{!��%��޺U�Ƥ�/^sc5��#�G����X�	A.�`�~���lYz���.}�~LNY�1�$�˙��,JE�9f�=��/�ġ9yւ�!��gn�>󃅀?�zj���K��?MU���a��Gnt���?��^��99 ��n}�V	�r���S���+�A�Y ��b��@˻�>F�dG���y#C�+U���QD^@��.�[,Gq �H^�k��P�����Jhd*7l�'ۺx7�NES����S��{�0f�ȿ��"{n[I��Sr9�XD��ߺ(��KzD��ؾڤz�R�ХM��0;_�K��͊�=Ya��#���
��Z9��RC��oq%��	�3� �>���:n�?0#��g���Dr�[�^-���X`��HS���̫���Lؗ,���l���I0���y�ɜ�!"��bk��/T)yP&̳��^Y���t�xJ���.��	�N�
�1�8���L���p��V�+o����� �'fm��W{���4�{?��{�o9��ll3r@�{����ۃ��* �A1	���=Y6�K�t=�D�ʱ���R����h��t\�8�7?�����5�k>�¾�xd�6��h�����hy��ol`-
#[���\�_cC�_a����!	�j���Z��aʊt�𤃜P��H>����j��	�6�6��/����
p����N��D��맏���-G�$Iw�1�(N�F
F��@P-��Ô��<&��ρNw��zB8M3=����<�irT��>������y+x��� H��$(x5Q?���e���>� n��ݕ�l���xe�^��&$glc�ysϴъD�1����ńh?��O�hO�ط(��C/~��я�@3�0pi�u��V�X�Z��ͭ��0v�ʕ�9�qI����������ŪVo7��(����ʻ!e�!��V|Y��ڽ����Ys�͋m�m�u����M�9Y9��R��h��Q�L��'���j�_�o*E�DQ;��%tp�'U��q	��Ⱥ�Pn���M8ٝ�O_����]�Գy/ �@^��&�������)O$�*G��i��J�.e����/\zv����u߲�)G�b�\-d����{����B�w�_�d�b�l���5�n���q��XS��Zd@�S,T%�y�~$$eIAU�>�ǁ��k{':���
�"���X^�x	�mNV�Zt>/�w�"/�$�3JTh5ghD-G�6E2�����uN`V-��/������厃�Y��"��9�_򐵅j���$��@��d���X�-pt'4T��g4�wS�)'�*@�Ne�K�������{���X��1/I�;��E�Oq��0K*�piQZ�c���5�0�F�UP�j+�p���������lq8D�F/d���էS��wqS�/oAm�k"� �Wr�5(�k��4*��������q��%ж8��Ύ)�Vomj�X���0f ?�+h���H��U��#���Z���7��1��� ���eY�h#`z��	"y��Y�'S��ˮ� ���͏<U<4�+l�^jO�\%v���LûA|K�*o/�0����D ��R�����v�@:��w����5���&�c���Wm?J�v��U����e*b-T�5`C���H�E���>܇S:���2	�g��D�5��$@����=�]*b���C��n��׈��Dl8W��I2q�-WA��9)��5x���H&[���\l*� IC_RQ��܃+o��l��kKLPx�����'���و�|�4�jV��:�v���p(9��;��_e�`M�;��!��M���Լ��)<ыE�j�3�p�'\���M� ��g�[�
C�+Y� n�b�[#��xO�T;�����VbHI�?.��zW�R�U�Ad��GG�[���kȗ<Q۬�^�[>���f{d��g���q�\�Ф\d��MEc�Y�;#�E���^r7���_�N��k��i31�+���ێ���z�k01��
u$����|�RVa���I0���$O�}�C��`6e�:������5N�6R�7vI������!���0�R��掷�B�J/6j^+�yYC�7��]>�m�g:^_{+�G�3�]��tPNt=LYJ9�pdrh�������Y�{9��Ѯ�'%�X;�!�J�+����X)��F+�1��+��F���Ȱ<h	y&L5� �k-�2����8�|�K �7b�{|�É�e,_�(ЇMC4�Rx��@۔`��
T�NS������Rh�t|�M=��h�AD�N� و����{�E���\x���Bƕ�aR�T���[{9���SlyA:�B���aB`�AQ��T����c5���I���ݗ�A2��q?�A
�y	��zR�yO>L(N�c�_J=.n ���ua<�tcaԧ�q��n�(�����Ɣ�ۅ�4<2=�Sm���Q�mY{�g�8*J����Fcp�Y��\��j8+nukZ����y����k���	/�V]/��(��mC�5=j���gxz� c7�S�g��H�y�B�X5�& ����,-�X����}�[60���Y��:8���1[Ȧ��+�H��Q�Z��˰��⹪��f�N���&�����������H��n0�->�����u�e��>�~'Q<��'@���Rq$���!/G�f��	A�N�울��{�t�#7��W��T�?�gk�V�	.�8��y�-}>b"e�"��ʓ�k�(qC�l��f�� 9Neb2#no�q��Ь��D�XvO�]kw�q`!�h�r����^)h�[N�:0qz�,焵�j42� ����!P�hw|�zkC[y5Ǐ�RP�@�9��́p	YՔ-j�F�{6\�?�\fye���B����S$�b�� v��K�W��B!f	��ر/ct�u��	��(�Rφ�y�KL:S��QV�N���6y(�p��Y �����)Up��tk�Q"Љ��iy?�搦��?�_�W�F}P*<M����-Sǝ�֢�H'�@@�5���e�v1��?�A�1d;{�K��}!��qj��������q0��y�9ڊ���x�����$�'�`%-�����(��wExoy�o�s5��Vhd�rY�T���a�dl�jO�[J��@I�_u�t_M��i��(�;.;x��!ѿ�\y�sȀ��(��c��\s��������ϱ7k��g�v���UXLWׇ�wd �vR�O,�'m���<D������g�;�	J��J��$Ҫ����w�T�eIv#��0�SZD�?=6�k�$萔D퐦ͽ�����|�'��]\��i�a��~0������t�+A��׹���)��'���Nй��; π[xB�A[uƨl��m�N�� �i��h
�����%��$כ �4O�i܈\m!A��}����9N�Hb�����')�(~+k����G8���҄Lʆ�%��OFu���B���a��b�V'We�?��t���=f�����P3�-��|Fr�T�����)ˆ�oρ� hv2�tV��
�c�Keu1�t��BB�̙|����!l[�J���cc]��吊��<�1��l�Q�ܒ���Zm�@��<��\�icZ�&���#�ʔ�wN7��O�*�M����P�4����%��9gS��N�v`��/*�E�	D� h'�0���1ڠ�9��N���C�Z�`{	��uڿ(C˽
B/{2�A���#rP�0��^�TZlՂ!vB�-p����%��$�Q��W��_�e��\5�rq7����1�J�������`��TvE��/��.BߓH\��w.�w�܅1���ouqz1�SחJy���~�6��S�(ֿ���^M���A,C� �\Y��^%3��� ��{E�u���g���ƈ�<H�(L�P&�G`��4f8����I|`�Ɉsc?�!����y��FC� �mN��S�Z+����u�<q���r�e���r~��7Q��O�
��&bT�4��3bZ\E�������b���D�Wo�S���L������F����툱����7'T�E��SUx�����H)����u좮q��J���t��2�T����+�B��>u}0�����[�c��1�yT�zT"�r�I	c���N I����S�"�n����k�S?
bs`	��f�D3�E����R`�hTqYN������Q<�;�Q��ɨi=�]��g���neЉ71�K�;7�3�#x�b8P2dN�����:+)$?Ļj�Iw,�N���A�5^h�&����ia������[�U�%�I�cS�N\$0G�l��5���qJ�"���)O���ז��so�t�f~+��
�o�� D���K�l�q?qsY�4A�Bh�t�����6���}KK�O9�V��?o��
���
�Q~�^d�ūLG_��p�q�D_	66��x;�wzщ>�tZ�V]��py�)�T�d05XM���寖���%�g��8y�n�0��Q������)�37�#��(�M�0A�B?�Y�WU�c>Q u��֕LS��a;���aA_	[���7�'��.�y(7i�f�v��� ��=�8"�ٚN���ޚ���'�/W�K�F��C�I���l�z��E���8��k��R��`���==�y�4a��ku:��?"�w;@�Z�0u����F-y���ZGA��c��L����(e�\Q1��b�e�pWb��w�X�f�I�N�����?����KA��~�l�����hq��p\�x	��\���d�Ȏ��v|4n�T��SRh�[�'�-d�h|����&!�Vou� 7���Y�.��0�G�#���:D�SB�9{"�RR��@��@�p���0o�5��Nl	_���A2�����@Ax�I��8l��m�Z��(� �������z�nG{�0>ٰ��ƣ��Ǖor� �O��x�/t*J��'���g(B[I�վ=����ŜwZ��Ê�>��D�'v/��,r�r~���N�6�F.�ֿ>Xl�At��ϰ��In�g��~Ě���z3q`��n�F#�	��M�?ǌ�v�dtz e�Pq7^dH�B��\9u��X߼P'�&��?xu�L)L��+.�'O>���B�4� 9ӂ[�Ť� ��غ�XU8�tῈ�#�!!
�VJ��s��� N�{XO�R\�����6�����\�n�t���?Rh���e��5(���B!���\]<(�u��&p4���~&AE���s�/�|��,�QWّ"-�y���*��I*J�=����>��vhi#�qF�2�౑y\���w4���|��"K*t�����?c���%�S���5xUng����}��oo���^i:UnV����+[Z��e�)�f�q�R���u�����z�+�Aa���J��qGl�P���
X����N{�v9*�9$\�t_�[�V`�"\����u�k�����Cf�M��՜敘4�֯)�8�]����6ټ$THQ�#����=_��}�H�*ͩJ��R�����]��!�$ͺ�B���ݤH� ��fn�7��`׬�y���X������!�EU�0H�E��4�p����I�E�"S���g�cw��@2̣5��<�x��k|�rXＺ��F��!����"J�Ԅ�hP#hJJo���V���A|ҩ���]���(��n"9��-&�ĥ5����#s�i��}8�Ō��O�N)\�D��ǞL^��tx5���bѝ�$r��Dӹ�|-�L�I՞w�5^H�T�2=)z�64vE-B:$�V�&�.?�kxE��k�̪����nt�0R�{�a/�{9q�����'��e�ڙX`@l���Az�ja�����ZIp�\��F��J=�
q�i���`=����xh'B%� �񵱊����$.h#�5�ҕiM�����3��3P8c}�k��bx����4dY�^Y>�9 ��~�)��찷��{p��z���r5'�7��M7����E5�vQ2+�/�Bq��ȫ�ķ�t�b�5U  �*,n9��!�q$�)@��D��7�L���T9�{�*�r��m��
/�Ƴ�ˎKIي��S0�$�ɠ.liN3T����~���|t8�UW������� ��E�j�:5��۪�!�"�֡Oϝ�d��4. �z4��Z~gT�P|'B�|�n7�w�}��~���(>QQjs�@��%i���F��B�Gi�{��.H��*}��Y�kh�#�>l���w�\�T����L��̮�^4�^9��ގ�,�S�?p6���8kjə%��o�:v)��"�Z��c���A�2]�=$�S��)��k�km�|1<_K��|Z=���0U-�dt��+l�E�*��9��X��������6�i�M7��d*h���JF���h��t8��Vf!�g�N) ��� ��7���s$<:�di����ʛ��'��0@�I:Rv�� ���z�GPh 2@�c|r��h,=�H�!o#u�_#O��� ���>�����	��s��b��g0)�h�{���옛�Cu�ԁQ���ŵ����'?�]�f�[��f��?߽��v�����=�%�{Rq�@��]�L�}����ͤ��~w�w'M%w1d��L~kk��K�� H�2�I�+xϒ�ZR{�Un:i���Da^oR[HC��sW����S�.6����O���޵��8zd�D:G�W�r�i�	�ĝ#Y�O3�i&�.ό�-_�n��[Uk��|�R7R��
�-�V�o�m? �A,�w)u=����WG�j��?7!N���R���-��:�qZ��(�|YS���+�j�B�]@u��MC��_9���H�.�:����j���W�<}vW~�ǪC�aw��<Տ�����+����B{s�GD�5�����@(��w�FM��=9��<ᛱ7���Lv��Sv�R�?�|�w�.�v�,.+?���Jd6 '��:�
�A�@����؏=M����Z����ļ��¾m���	q����둙��.`|pտT��3�B��N	�q�^�����Z�Y�����M���pu�,�%�I�}¯84��O�����r�
p��~^�=�e��높߱^�dX���@�C�����i��'�c3�v5�35z�wQ;��zvI�;+�Ѹ�,B�J����U~q�r�~�H������g� ����ZkI��F\���d���;z��<�5%<3^u�|�Q�2�}�p ��~�-A�������̊�gM�Trn���)��m�T�P+g�V[,p��45�J�'�W�C�W/��.�4:ؓ�J�u�]�Q�����@�1묶VXkԚwM���>�aq��A^6ʠ�h���HS8��QR&��jE|�;&-�5yrڕ�?]�J��@״D$�0�/@�+
��	µ�,��1�C| ��KiK�\�����e�P�B���V�	��w��j]�IJ1j�%%����;��"|5ж�k�g����0�.�دg�R�n4x�D�{@�k�,{��{T�v��M����}��-�E\�7L�ܼNީ�fC����u��q
֧D�u9}�d�g �,�!���gcRQU!d_�[2	�М��1���61x��Qd�an���p4�Ĥ�\Sn�{nyV�qy
�|IkGCl��U]x͖���/a.�'w7 ��Al��a#gel��a�@ޚ��
�}(h�)�Ť�,�,wuD��V�X8��V�B�	VC�p��1�ɋ���4#QԘU����}����%]F|�,G�ԍW��d�F��b���e\GC~? ��I�j�1s�!�\����|�_�s�4��iA�ߤ�
��V�b��޽\]ҿX�U�nI�
0��;x�Q� �������#�;�*���5��n�8�u��f��S�?���C��C&+d�Yp�C���c}�)�rY �P��@�4�ewq;�ӆ�����/@fj�Y�E�Q��ʅ&v�T �;:�8~�������|��Ρ��J��$te��H������_b�TVZV����ַ����f�n�P6Ё^�|NSj{%��jF�� >��w/�*d�~.��v	z%ɞ�lr&���[A
p��fO^ʞ:�1�)��{nO�v,v�G�i��MH|��x���F�=��nE�����u���u�,���K'���%}�����\�l�۲bC�z�e��r�9H^9
�@�|�P�,�;@�e���8�0��Њ�iZs���Jv"JT9��~u7r�/�N6omT����(���U�C �;S�ء.N	0Jx�Ί1�'�f��Ϳ!���
�L�T��{��r<�#q�P�5Wz��jpN���*�9.����R�xA�����G�Q�����z�tf�M�����Ǽ
Y��ǻ�"��aP�����?"6���G~)�r]�J���Y���m�N�6����o}�\���:�ϛ�:E��:v�q�A�8)�d�!i�A%ƯH�,y���b��Gc�6���.�zR�T�L�'o3����?[k�u�ũ!~����g�/!�A�m�ݾ��� �Gcb�נ\j�����Z��'�Ju�OLf�_3!)������S��iW�[�ݗV)�W�*��H{j������O�UE���#��Pc�3 ��7>�^��M!`���S��$�/|h��d?8~�.���?�l�Bf��S���e֣l���W�6���T���X���1���-=+�K�Z�d��B���wO�C�-m�������!�{r�tQ���g���B!G5W�� G3�l����/�v2#p��z���_/p`?`��XC��\ǀ���4����]��wC���ɜ���*��D��m�֮ЮĚ�I�Q������mǟ��@:�j�By�m�0��DZ+S�WL����IT��xx\_Tkw�����^iН�+M�ܵ(:$]#	��!�,	��d|���M6���1�!�Q��uYI0�����.��8CE�~@�Ű�Y�=�F�%�h!M��|�C�M�O�Q�w�^%1FA��q#��T��Ja�1GBmC�G��_����Y�B�or�$춓q&�=�V�����K(o{�z��E�g^e�E:����S@TmD�N]Z2]f#���?F]���~�V#�\�BxJav��]��D���[Kf��q��
�xu����3\M�!���ɜ��sI�(�x�'�y��v�� �*���^�țb塠�#�γQO��2�ŘC����w ~��E�UQ|�V�*C�!KGB��*}�)�F:$�L �$7 t��X�uZ��s-m����)Y���Q�J���Q���<L4fSy����$��\RF���<�,1߆A�G��g�/Gp"|ƒ�հ{��i��ߏ-1��a}��zmԪ�ˌ�e)���%�]ګv�`"��ϓ�|�޳���xR���1��g� ��KXQ����I`�;�z�*UT��߽�9��L��3 c�*_�N������Q�����.BI����M�q�m��11�����^�Wt�>��f�c-!�*�W)��8��z���%���l;S�7&�/Х}0�7O�p�j�/M��GI��x�8�>K����H���\!{<-�w7�R�q:���a��g��^�G��j�轊|n:T�/��:@�;E�=�\]���b��/�u�M����lW��q�y��W��������qb��>��Yf�4�qhT���{�~��d�K�ԇ_�}�.$��ߩ����=���g!���5U�zufd�p�p��mݔ>����X���[WOa����#�!^U�Y�z��|�j)�S�
���m>�l&��'������QXRޘ��{��;�[�8?͵xu���(�Q���mGxn.��j����E�~XfW?Y�]��%�B,�c��ױi�L��z��&*Qh� �Q�O�"�^A�M����%�wk7�\��-��T��*F\Oܼ�1��aƢ��\��\�^i���ػC4��6��}��%b�1������x����8��B&�΍反7�� ��+�V��zsj�D(�F#�}��ti	��R���H�љ��^�Rt�C�������BU��OԂ���@ݜ 9�%����c��@	�E�~�`+�Fȅŧ)6{+�yG/��%X�J�Ԕ$�B� dS��Y�PM�,�b1�*�,Zw̽�K;��?	�⻇ʬ���ƻh��sǄ?������?�V��9���4��ۮ<�-#e��t�c�r�m�m��l��>^�m�ߦD������^W���%�Ƨ��4>ך�^�|{�׎�d��@@� �=z#�1������/���Fl-v�=0�ZG���|�cҞoJ<b�}��˿���E�X¡�eH��r#m�oO��Y��B7�̯�`��&�U�5�c�Upc�u�Ĭ�R�{�vui'�yE�pꙍ�?=-��8�D7�b(�*vw���\q.��xlq����:	����-��R���`�^B�t�T:-t�+&��|�ȯ{�����7�W�D��W�v���HsQ;�S�3�Q�ʍ@�m�i��@�BCyVY��Бp��5UIa�{t)�v@v<ʋ{�Z��WH�8tQƫ��*(�sG���:�tUPB*��X��4q�w��澒�h7O��!��u��XY��S����������`��v�u�Y5<%�僣��tL����7"�+ӖAo��=��;��7���/T-_@O��=��)C9�w]٥����/��{ 3�yo�NH�W	;U,	Z���U�К�$��"}��5ܫ5 ��K;.���c�X(U,_<��N�[�����Z�j�uM y���^����Sfc��ĵ#��nL.�t�����.u�Jl�y���O�S�z�!�P�w �)j�_"�Z�����1*A@�R��z�`�q�g���"�sڤ��C���� �J�_��!��Ђ���,� �G�8�or��� �r��qP�Eh9�?�r�zq����q��Z��'���t�z˷ŕ�P�Ж���<��
v]��؝�A��̆n���̥Pr�f��he�C����RS�)��D�R~�F-'_j����ZD�,-��6��r�Տa������윾(�j�H�����#L���klBb��%����-wL�m� �e��w��at8ƑZ赣0<+h0�,:p��N���N���W:`.�n�BO�(��;S��gk�ٙ�E�t�[TL��_�Ϸ]֔&��1ݱ��Ǉ�.������~��K쐎��sSٕ>�s:�$5	�)�Md�=�gǆ�����CՈ����#4�P＇��$C��,�;T&*�]�Y���,�qs��$�V%WX=�^n-��A�:�4\�3ݟ�V9:�s�
�2#��C騖���y ���5��4�~;�~���UKN���$SOr��Y�?Z�"�Ū�-̲���n�E��6LB~�JVr1��.��K��&1����x����d�in�ͮ1��ԁ_A<�)V�޻DC���cKA����.\J���,�IV�[y�die�J>�y\y���\\�dZ�m4d�Rr���0S�����|��|k"�p���OIѴ�u�e#��%�(�����w\FQ�����?_>`8^�K��h���/aY}��"M�B��u��Z�D�.����&iRb�d����ݝ�Z��j�~]�uM�w�zL�*g+2���S�H�V2��Z�'R���������O$�([�Q�����xY3�޺���t_Ц�Jm8��;��^6�z T���+d���K��D"T��9B��D�p@��'>19��aT���<w�؆�`��3�N�:iGyGgؖe��_y�kz�����U҂�+D��\'ͮ���$��f�� 议:��ʂ��lPM�?/Հ�$��i�	xK���F�����UZݮ�j�h�=���v�'R�-�������n֦GI�� n-�3��2� Si�C��*�1�a^�U@��� ̓�4#��\GOB���U���������	�U�������&8Ճ�)aFrh��F*o ��Y*WVn���S���Ǘ��ww
�x�-+(�0:��UCN�Qec�"�F����uN����52�;vCa>~WXv���je*"\7+��]/�wo���uu��┍�I �ZiQ�=�3+cs'}8�}�P��Bh���[�/:��|����[����5�:K7�֡QG$��Ed\e�9͂P�ވ����Q�����]bY5�` �J�����z��G9H`�'�^N�z�5<�ȐS�>N�k�K�X�wε���p��;�D_�3��~�ش��" ��B�H�sc7g���/*���<�̂�K!�<K�^~��t�*͞�|�����L?N�.��ۋ�A�i5�`��L|���s�CU)������n!�6TY)W�(�Ã	�엦�G�� 4+�"z�jx����VI7M���L���􍃖xzOKe�9{�mL��1l�.X��UR&�$$[�]��\	T�m/��Q��8�Pw��h�[���$0��'��,��9?�l�+�gHKa�S�.������d�����Ew��pz��d��ә�s����'֋qdK��!��t�5�}VGPG�׺��;���Z��X���A 9�Ɍ�2���3n�(&�[I� ���}#�>���=(�1�v�{\�������wP}����#��K%�wk�ccb��TOI=��4��ƿl# �gi"�ڤ�Ҫf�
�r��&R0�m4��Z��If��>�k}�ҙӜ�!i9J%&��4��3٘L��]w�G�:�=�0��d(�`)�x�a�+K��9~p=�������$�'+`�����@����� ��)0ɤD�h��0�3XΎ0U�2�V��\CFߏ�h|����I�n�3؃��u�"��j�o#v��<5X	�4�D��:�(��}�߻��6�X��~�N�!4�H>�$6�@o�L�/j^\������(�(�m�Q�L�F�S��Z�V�^;A���O�䋘�!�<��.���u�˝�qgm97?��� "�b����t`�V7�)��`A>�����rFgG��c����fZI�G�|��[K�sp���m��G�T���J�5c�;x9�;Xˠ,�z�)q���ɤẆ\�R������`M`��6ya)�u����$�0�����}��z�\=�i5=h��6.`���&����N�?	a
F�4�u�e��Հ��+v!�4�x��y�F#�4�Q���r@�i��Wb�B�u߇��}�[�^$��2�̆�I4Rm%��3��Ҡ�VW��G�������'/F-}�	\�l>����z��c$�T�&��8�¼��3���gnAn�� �$�>����$@�w�$��^e�.�󝭹���L_������� ����r�c�.�(Ͻ�*����Y�	�p�}��T���թ�Fz*C�<�����ˮ�k+�?��l/�I�i�'"�ʦv� `oE�&/�/c��o1�Rf�(i/��0��Ih6�� ���o�C\�M.����b�rⓛ��e�]�gUH?�nFKa�U|操j���̳�\��-nS8�%?i�ߔ���v�f��N>c����]|���+Rs�H�O�O:�#���A"5���K����F�x2�����7�K��l=}�o��xN�����:�y�J�Z9�D�@�&�������sm֞i���<2��\g9(�*���݄���s���}<�&=�9=�[�Be7f:)<12���s{F�㣍�^W(m��0d�x�73�T)�5��=�j�*ڇ������_W�����餆���^`�i=$�	�st���- ��>1��¤��h��~0���)9�����d~|�<j�z��/Z��E�P�gPuLlZ[l-]줋4S.���&����U��me���FW�.�̿��*�>iu��O2����M9�k�}��r؏�b��p�%hBb)��0Q F^��熏�M��O�@p���E�i�N�sx��� ����G50��ﵕ&���#��N�Ҟ��{��ʁ5e�&%�	e�[�k�P a�����h�����w�Zr3�a�V;.l�i�7�Cɽ����B}���Gmu�p����I��L�E���;$3����>~%z�s>�6!�^�R|��+]<b�uT����(o3�oaae��Ѯ�T/���q�v�)�M>ӽD׻ϳ2�O�˱��S.V�poS�ts�S ��{�ޑz�c\�c6M�}�\�c+�������GI�� j�`<�~�
bט�Q-�~x0���=F��mR%��=P8{����.ߓ\ N��dm,� !����[�����	";*��K#�@"�O�h�]h�
��N����=u��N ;�Y2j���S �&���(��CUN@��re@R��e&��A2�&��5�!Qθ�ٲd(�ND��+���L�`C��d�?��"��!��*Vw{���$�j���t� Z\1#3K׾�g@�ௌ�����[�g�z�\�h,[T*v<b*h�噐ڈ:k���'L��
�����  Uh)u���f�?�5�\��O�3�Gg?��o�|������as�C�CF�jn$�rIU��@�Gyc��:W"G�E|�̇<�=��}#V��(߃r�~�L�~,d8B����`��)8���	�h9��R��1�ߚ
�����w�A��|�b�Z-N��[q��a�%�f����������w9�����1�h��4b�Dq�&�����t͡(�~�:�B���}��J��f�DAL�O�f�G9s[�?nTD5�Y�J�vu h��ٍg$Հޱ��䄉l�e-�lxf��A�-�/���1�1��My���"��TG������(�t���I���p���jx'��hQ^3nm��ba\Cq��@)u|p�}�J�P�#�NR���UpFȄdC>�"pt��1��!_���N���_ǭ���DBAk�"�/�Ǚ����tEv��~_o/X�A�Z�"AF��5i���q��sl�r��3��i8�9�J�_�apK�l_Z�\�����)5�}ď�Qei~��xLb+ū�������_�B�8b�^y���۠0F�˴T�ч��IGB6�p\et^{���.=Z��M7���t5>�	����4oh�4pv��b�1��+��G�"7G���Q��f�BKա����퓨�і,t/I�Wv5��X;��籛�/�0�g�;o�Җ2���ho��>�����m�F�]oځ��U���%y��l1�>f�_'7�hgB�⼜s3}�����IJ��q7P�J�.���J���+��h�!�DK�glxi&��F���=_�3�ǟ���91j��<���>����zŰՠd�{^��}�ou��~��ٶN/|��j?	�y�-�s���Pi���z��J�	�q`}]��m�~�ug���V��V�$ca��70���~�(5 F�`-���W��co��HدÐ�3Ҳ����h����)�G������~�F�ɟ��d�A��H������9	9^��P���r>��H�퍡U�vϺ�.k�T�ǠcY��٧�R*��.�o�3�5#p�}Wz�~��� p�ߐd�ΊJ7{�O\q�0���wZH��i�"C�~��+��FXb��2��')�8 �4�DQ�&��Ǥ^]�K�:�k�6`��5��\�a����s��#ar h�g���^L��Fu����6U	�ms��+}��3��p�u��:����]��jAP�d׋ʱ�G�h����W�4րgN�f�-�Q�ws#q�z�����ɬxN��޺8�ϝ9��fC��l���]�o�ƕ�!sU,6�X���Y*IGFO������s5�I��5-�{�pbdH�@��1h�/e(uں�M�W�b}?D0h���5�m0�t*O�J*�.(���z���b�70�[9�dH���K(w+�][M��Z�`�(?Dw��ܒ�V��`�-tv����6b���?���NVD0j �\�J�"��#|����6i�p^mc��HL�������Uc	�y����ɩz�oF?V�����G9Un��B@�6�[_�w��f�
m6�Lh�	��n7� )K�@v��.��X�$jh-F���PW��֗1����ȑ������
ؔMŠ�$�(�n]�k"I2���G'6M����?���l*�o�ؕ��p����%�2'���{�p��u�&������Z�I_'|XI�U��X�4�)�ꑂ�!�F�$~�69a�Q)M�#F�E��Q���湠�Ƣ������+S�Π�#�N!�;��rH���u���}S��H�������9�1<A�>l6B^k�Pl���7Eފ��h�Y�Ʌ���^�*�L8$�oWS_��^��t��Ş7'���5�}�Ha�!Q�����'͎�.	�1�`���R߷����vlQH�_�'�c; �����Gx�������Ao03�g�md��k���P`�� �\͏]�����۳�+�ѠJG��*��L=���%��>�'߰���\�?i>W]]�>��PB�O�8�A�Yv3�a�gum�
|ER�u�dW��*(BP��(o�V�=f��S�V�(6��C��_$�ש��_"=���Q[����U�/�]��,��£1��o���wGo�A��x�m�?B�gss�80T��8&�<!.$���_�JZJ@�ⷕ��K�缔�;aIv'g�}�w�VI!;{|ݎ�N�g���D�j����+i%~N@
�g=��z�ҨbЙW�-';�͈ܽ�dZ2%�fX�(~�����0^̖��:���2e�d��7w�At��0�K�=�3T��sۋC����7�
Ga�I`�+q}����$�;��Ŏã�`���N�H��)i�4
E
��y��'w˫V�mO�v'�&=�qwitr|�N)�(���Gٴ��0�f�5Q�z�L̊磛Y��M�G�s�,�a�&m#ZϹ���R��a R��/��+_+Ɍ��rk�w��U�&�\�V��Ȅ�g���4�EZ��c�v���;Wu	��i�����C��UX�@�A�M֎&���L_�~�բ�s[�m���bP&�tJ��g����?���o����k���b��,҃�\���TI�l��.i������ ����i��}�I����q�nLFsIB�ZN�˦Txʞ&��~�deDp8������}������d	���Ǡ��4�B���ZV�KG��� l$��,�]�����X�K�?�D���o߳@8�8��<!k���I�#�E=!�d�ϵ'M��g��*nL�11jAI	Z�.�ri���)�Õ�!����T��<��1ݘ�!aX�w�q��žy�SR�n����X9;4�b��`��Ҝ�����iW>t��~���3��w&����@�@�V�l/�oʁ�	9ks�N�w����Q�[�l4��ە��
�/�`�*ہ��j�tP����.^Hb�j�$fט5|nM�b���l�l!i��h���u�+�͋�t�j[����4�Ny�����������No��Gf!�d�����ܚ/ZcC2����������/
Q�ǟA|Z,$
̑�B�Ť��!kP�����_�m��������Mg`��@��zÿ�`��>��QU<�A��zZ������a���X�+�;�=���H�%�C�J�G^UuR���kû|R�7'�~/���D*%%����*8��L޺?�;-�CE׈&}�h�j��}����=rظ��\���<�u���!����U�p���fᏼ ��� �wkL�B�l?�SD���x�We�UN\�Ƭg`����K�;�
�?��89y� >ךH��
�7��@%H�k=�胝�ïE�?�!�2��<�.#��$#�%���-�*~�\�ߴ��WMf��ՏN'@z��w��~�a�>䇽4t���.e= ӭ?��.��W��=�>=�HW/'cvx�1����(P�9pz>;�ε�J@&)H��n=X:@�?�>��\�]��P�����z!��+S9]m�$d�.|�x���T��K��K�G�<=|�3<��OuKBLj.>�N��$$[��M�F�B�a�3.��_��߸��)X��^j� ��I�fј�χ�f$C��� �dK2���Cs��x1��`w�P�`��o]c���"g��9��l�e���x9e�f��ω�;��v�W����1n�)̉�
k�B���CY�<˾+�\�^8�P	�乶[�*>T(3�Ո4Ju�������O�,�0~.C@�I���՘��ٵ�@�	_�M�hYҌ��� �̲R��t�)P��yX�a�u�5��<��f���r���*T�&-�	w*��sLX��n��ӣ��$P���]��8#������N��ʇT�3����ƑC_/�f��3.Xĵ��̑v�7��B1D�i���n}�@d�	����JÆ��M;�YQ�F�xX���0�׿.���a���Wl2�z��~i՟�8�R(�cl�3�ߜ�喇)Љ���&�G<�[c >Y8Jq�V��Z�4<���5�2�N"�	�rI��x/]g����Aܳ@��$@�gs�b�J5��oqN��"��zn�ɨ�K%8�J�C��C���&�Q�w�oLNFbe��:B%s| S�JY�d�`�R#�N�B����d���,�L�1:2�a�C��Fl�n'������`��zE�tx\���h�%��L���)��1�(B�1�[FwF_�>�b˺�酞���,<�9ӄ�/˥jzW�D�s��<q {��6D��.�w7��qJ������'D��P�[*-�]�w�0dه�F�:�1ꏜ�=sd��n��0�S�%�V\���u�s�=.t/���9���EYg��d�b���s�^
�_o(��)��vg�R������*��q_+*;�����&�H�)��B�$�"�����cЂ6�����Z�x�h��&�F�������V2�j]�`���Lz��8l�I�*.���
�)f���p�d�ω�qZ}X��/7����م�a���q�r�!`��t�ݹsz����2�b�*�cZg[(G�Ť�vs���9t�IP���Ե�p�����%4�WaCL�
��ːN$^�oI�����'6��2{����u��p��d�D�h��g����;��&��3$�E쁰��T"�*�y�3��цrK��eN�qn;|��Qqg�� ��ߣ 8�����cR����f�[f��2�֭f�1l?}UFZ'#q
l���ϥ��\(�xar�v������2��)� ����`�C7r��X�?��JgC���/X�x�zE�u߀n���9 *�&'�y�3���c>w�D�ڮa,����?��L��\$u����SY��B�0�6LnO���zrx�1�`��`W"�Ee�*���3�©I�@( ]�%��e�u��ȝ~E�P�J��^������7�PP(DDS�uc�d5 4� 5�e�*åG��vNP��:�@*�9�u�OU.@8�*N�觴Wn��.�����r޻�ܛh֩�]���S�Tki��7U���p=C�X�_�D��4m<���k�%!jE0�RV����⿤0��p�dr83��= ��˽ɔ��<���N�*%�D�dVm!�P'�6�`ȹl&kF���e]���p5-ʏ�� G7� vb�DI��׮^����p��xf(p��c���#�x�M᚟j�L�!N��ꀙ�4�5��Km�k�g�m��~-��O<������7�՗����h��ˮ�ʼ��}���� �f���J����+���,�(p���9M����fb;�Y8�.l+��+�T��/�[k\k��;�[��Q�M!�=����N�'�bOWD�'f��V8���<!R��\�|T�Y��:�(�{Dz�b�(9Q{W��n��2:=��;������>�Q�<+�
�˱�K]s �mGb-h6|�X���gEi��ĶcK�
�n�����+�
x2�� �ԟ;��̃�*N��2�v��z�[�J�O`����;����ŬW��).���2�x�a��W�����^�ݓ���I�X	t����Eҹ;:�~�����K�*巓���qZ�i:��Eݰd��x��$��E]�FndkBȊ{8�s�l�5�����H���p��?�D��ov|س ob{����D������mSv�j/c�]m�S9"o\m��ʍd�l�p؄���c���~�y/��^��ܐ0����SlQ�H�CiʀN����_xUT��#�ve����%^}�_=�� ��>���*ֈ}{�W"��DG[�xn�:eb�'�a}<+�qctO4l3�� �K$h����(OV�"B3��dӱro��ϣ�\5Tf5xͷ��2�Aej�,{l!�S�g��ͱV��ҹ��o�L�3oH����7� i���oPO�T�?s�6S�����O�3'��X���f����,r�B1Ŀx��J��-��酠F'��׸�۴�
�Dt��cg�{�B��l���W�����4�'�1��&��5y������笩�à�r�z0�b$}[���)���κ�&� ��z[ѩ1�5�+�u?Ͱ�u7R�B�j�K1�g�Pd����us��2gߋ{D9�~>�[�3�M%+C*������յo�
����02��4��5kp��F��.�jtvn|Cѷ=P��#h�|{G$�\�jWk�EY_c�7� #B,���-�}ʾA���^%e*���xդ��"y�&w�]y���V�B�����n;HCX�0��#f�ƋƖy��y�Y5b��,���$�W
���E��,����F�2lͦE�E?�/�=yϊ|x�����D������	)[�ߘkP�}��g����3l7�qf
�J``�����sɗ���Ԉ� �A�/�оD�O�b��D4_ӽ�хv�0�D�X�Gf���|�L����D���a�D�����8�G��+���
IL��MGET$s�1�PL>B�h.����(���n�,�LLj��M��ܭ��[0k��!��<�tYz7C@��S�1Z �\j-I���y��_��%9��e{������4$�� y���	]�a7"�^xط��w +�/)�sd�s���j�h��jƶcT�:okǋ$��ɬ�� G�-�I��B���c�-CJpe�wU3&�f�Ⱦ/�9����ȕH�4�-�oc���O}������9��w�v.�����eJ]����p��	~�R|_L��77]ف<X�/cs�}���MA�V�C1�G�Br��9���l&V� �1<w�������95���x7z�(��;,�pHb vj��֡���ɫ,�/�	��)<l�s�y�xVMc0��s/q�VCY�bw�Ӟ=�'Z���C�'�u�K����?jl�7�:��DFR���	�Xk�oIlH��D��\j��~��W�ׂ+t����>�}5�LkO[�
J�v¼�DM�]J�K1����W��I���w�}��PJ�׏����-������&��ݽk�M6ɀ��>ۗo���/?�z���cwԊ�6o�R����X�T�x�)"�2�Y�5�pz��qP�۟E�2��aB��qyQ�љE�CC���9�8Ƣ ��\��Y��n��G�_G��@�؂��N�{Nn Dc��K*D��t�(w_�����/DR�2��|�`k#�D$��E���z%@ˈ9H�nJ�W���L�|�Ƥ��DO����Lk_�8݈�C�r㋄���gfzy�'B�[�$��s1�Vy�ʝ��B@��m�Q5����-��$�^�Z�Z���p�\�w��g�R������F,�KV0���
w��3��~���-�(W\��ר�l{&�^��#ă}z�+�9��O9l��$bW�%]wǢ ���Iȅ,�|F�G��
�3�W&nJ�k��Xd�'���d��R��R�W).ݝe��9|ez*�{ڤ��yh�L<l�([.�&ܲ(Et!F4O���>|x�Z��������{��N�����xF�B]�LFM��I�l^] ����H'ez;�n�3��J�ф��<��/�LH5�,�5:���P�G*��m�+��H��CNG��I��
���T�Ƣ�y�].�i��v���jL���M��WC���%��7�B�=M����ikXY��B5��������&�]��+B�ۻ��!0ңDJ*&�BjY�1Q��o#�J`Λ�?v�Q���RuLx�kA^�����E����Ҭ�4�"Uo�.�lL9-&31�t�*��{�7k�~���&'�]�(��d��\X(2ߥ]�Go/���:Y4-���?O%/17����|�3�0���XD���MdǶ{��֢I��K��:	<�U�KW?�?�Ӻ�B��rV`~-�$gk���9������6G��HL�Y[���,ڗ[sR���g7�'��Ei|M�@���|�0!|���oU�Q#4Mʋ�?,��@#�t�b/�<��g�tŔ֢�����yZ؝�����>����~V�3u��ΰ2r�u�}������9�����\D\�R̖-?卂Gs�9����<�ωd|]���^-ë_�4�Tc7]֗"�nDly�7��z�կ�4s@O���X-ۂ�Z��HWS����t����/�����3'e�ݒ�lKo�,rt��������qN�&�-�ߘxm�Ǭ��J
5H�̆��_�g�E�1q@�vq^+ΰ�����1��X�M\>�ϳ՟�T�[J ��R�!^}����~>�c=ܩ�s��]���w1h-�+�5hp��� �T���w�����=3�q262��-�
��*��	$��O�L2��;���@=m#�:�2ʂG��b�Ձ��*��������Fm��Ԕ���k�'�ZH�d����[�	v�N�ζ�*�Ho���Alj���H}�Fj��){I6� �8��3.?��zV�Vm
`�a��N��!��eWA�3[��?�t�Q���ͩrì�0���:�m��I(qy�e�C���{D��}�ӄ�R�R��-��-h���1��z����8��a��?��H�"M�"L�3�R3~����r�ۥ���&G���i��M�lC��mI�%��8.{<���>s?*z��k��[�Y�uT;�T8���$�ɰB��	����n�]v}EV6_fS��)��D�,[Ǳ��,�L��3O�*]����.��M���-�UW�]F��xr�V�F��#n�x�F�Ct���t�`���!]852>-�pd�w�Z�bE�,M̷HISKQ�n2J��]B5F��2,~z�r#(Ó�Q�4y{�� �|��s���Q�Ef���&sB7�	?���Mʷ����2DES���Bu���ۨ8l����c���qBƍo����m����^�5B%�ĭ��,�s~JESބ���`s$��I9�퇢a��	�O"Fu���e���ӕ:�d���� X��t(�J��e�zW�+��;:��ޅ��ud3�7yaO\y_}}&a)	�%�[�e�% ���:B�ʕcX�t���Ny�u��w9UsNm��0I�
��C���  B�r� ��c���g�_T��ޣ�S�z�Ʊ�O��aQ��uy��z{V�[�
��~�
`��������3A��KlO]Z�1_�5�KäW\Fp庬&]� Ǚ�Fx�]s$���\}���6d�mw�[v�KP1�7<T4���Ȳ�b����YH۱�a5�H�VA��T[\�E녾5�)2�l$ׇ��\/�[�lp5���vX��b 3���G���M�>3�Ko�l�������tU뜃'��ħ�}Sx�Mg����q~�`��SX�]�K�s�:QZ �N��C�L��K�K6��7��;4��/�Y�A"V5s[��%��n�Tk5nM��)H/��:z�'F�з���(쵟�<�SY�	�u���k$��ؚ�k+j�#}�{Îo��X^�l�^-�s�`l��S]5�x��?��ZF� L�}�[��m��j*�y��1a�����mmrx�{����h8H&D���;�m�`ui�$F�Rᗱ��_�f���Q���jf��P����t�C��Z%�z�*O��ϼ.�g��
'ء�N�Z�� �ƒ����}^I�I���P��o~i�^9zwT�����axFP�͗;���7�)��#���h���N������a�Tw��$}M^!G�M� ��T@b�X����=#��E�9w�Vf�����Ɠ�%��~��S7�;�F6Q#'����n+�h1��h�6���3�Lm�������"!�N��_*)��6>�������Ss�H�  ��Q��RvGp��k�G�YE��>��O��/�I�#�E?#��r?��3G""�&F]]Bf��7X	��j��I�W1aJ�����Z�F�)<���)���&��0���r�]ʪ�q�MtX�E��36�����'�X�(ُ���: AǶ1q��T�W�(*6�)�Y�a�:=����ߩB��ް�a[�Y�a��9.O��/i��
��H��7��j�$!�%Sbj����*w��B���~�?����N���*��!���Xb�5�x�o�EQ������8�괲�8��Vΰ�B�-IƷ�D|_����u_��;u8����H��ӷcN�~���1��I��C���_M�ʏL2Z�~���o����e�%.V��������b�����`��3\����AR�^Sn�}�Խ��o���tU�œ6n����#K$6TJXy
��%��ff��XX/���@9������E9�����
2�i��NBG�|L�����pԹ��q�D�h���"��������ՓG�}_b�$
gn緽�p��:M�V�%�ˁ��_�74�k�����s%����2��G\�aU�ǣ{��x���7�E�70I�2��0�6�I5���uf��� ����]�d9�5�����#d�-�n�Ғ�&,T֕$5�X����/Sc�	g3b"B��E%<�W�s�y�@[�N��?'/�V�4��r�̼G��@�	����(�]��Z�w�?M��J���6U.��U�$.�&x���΃�x�;Sޥ�w���`� Ho3�Q2�n&�85����<���ai;E6Ւ��)�p�$7YWP���%5��1禷��Vס��Z=-"���xM�7%�`/����B?���A��1���������dKwSdV�w�^�g�q&����L/���T�f[�u��S��7";���h�B���� a`c���������m,�Ɲf�ehq1FL�8���(@�ljЗ�؋LA[u�߻��Ze�'�Y�SAOo|��6����pڤ#����#�I��L%�|u�a��#�t����#�(�D��2?uܹ���u��8):�Onqg���f{�X���������y̬M>G���F_�Eԁ=�@ʞ�I15M,0�����L�"�J�lg����]�6x�"<G��(Kt�"��
���z3���*h�p�W��	�H6nT%v�,\�B��Y4Zv�Һdn�a%���>�ɩy�zˀk��q���F�A���%P4;�`]�v[U�z�"cNڊ0�l��{0 �8J�]:��M{����s�����U�ɵ2��!cMMK��O7�� pyDwU�,�E�3PV	-�@���))��`.�������S�Z��F�"0;3u! �Ni�5Xa~^Gq�C���5�w`��
)PX�u|������ 4�i�ɴ�-������,�x�Mdc�����t>{��]�!_������˒Ô��3i��K2�M�E8�i`5��`^���1R� x�g^�c6zo�5���F̾B�-��G��FzC�E"��2.m�joF�0�';�5ǅ����ːH��;�[�,su����xG�I��Z4Z	�x�`��+�^��|C����ń���<Rd駲��g�EN�e�_V���@�e��.��|�a�6ZR�=+jv�:������h�Az�D<Xȷ�e���ʼ�m���k]�Qg?f��k�^KƓI�xr&�;]�G1�ZE�#����
�ۀ�7bg�������g��X��g�aA�&��E�|_Ҁ߱&4 �	���‷�bUf�T����fMQѸ��x���s�Q(UV�Sx��8ֹ���{T�Wg������9F Y�>�qӏ[�<B��>�Y{��;E{����޼����bv'�����QІCa�ȥ-Ʌ6~�Iͯ�MN�U�g}5�~RJ�E���w��h��9�L�Un��կ�7i�A^��W˭/~&��#Kf/;e`̀ޔ⚂�Kd^&V
F���qj;�X߿�I����x\BT��L5h�sE�`:��inL`cGxBLEa�s���{uE��t���v�R./�-m�V;"��4�a����~��CeǓ_>��>�7�(���U@R�εv����2.�j�*�֮>I<�Ɣ	��(?8ۿ��Z�qQ�ԝP6����!7��X>ʁlHEh��Ͻ��Q�X%�vxC2*1��zߘ�y�\�M�^2U?������C[��X)*�޽`����2:��k�4��}] l������� %@Gd������SO}u�<+�FMg�?R�jb�-
���6D���BvU��!���0��)��hw����uo�柝������ˎص���sAL�`�ݰ}�Utt�\+ jL��9*a��'��#'F��n��0�&mq*iT�\����X*�	EB����ޔ�5��$ҏjz�b|���1H �* 6C��=�mp�fG����L{g�=P�O��s�b��U�𑓜"�6���LB�2��t 1ъJ;�{���_mKXA�շp1���ˤ�}r�����#�5�ž��`>���&��Π�Y��;�E�T���8n&]X���&��j1��q���Ñ<ɟ���Sj��ԏ	m,MCFe��י{1��6%�U�o=S��G�V��6��`����E� .D��wdS�b�\+�꜁�V)㿰�s�va\pL�[.�q(�������f'��VQ���E���$ҍt7�v�Bs��bpe]�|t#�K�U6���Ӧ�m�r���p�{-/�ߒ%ӏ>Zs�W���w�hK�E�Vӹ)]L��(�*��K��Poc]��id�����Ύ�׫`�s1���U̶�vx .��@�rw?����S�mY�ow�3m����l�|���q�@��.֌$���� E6/e7�9V(������`ӂv���	�m�ji�g�e"��۟'��hҔ�Z��1C�^�r)��� 6�3v�D<7\sq_=$hӊ�
"m i�YEdN��& ���3�U�7��
2�)#7C6���ΞW�\}�%��{Sj���e��ٿ���!'*#З���F���������j�n<U��RTʜqUy���cr������-)4ИM2�2y���Y/�b>��-��yv�_�A+T���6�ͮ e��m��54�9��q`�A��p���"��'��n��$D�&��`��)(p��;0��!عx���Y|[3�ql�<��/i���?bPwY#�	�c����6�2�R^a��V�e5*Xl���O���9�DS3���[_�vy�5Q4����B\/�~�`��u&�F�iJ�K���L۰����E'}Gl��Z���L�o��8[�ޚ�f�:�O:�~�m���"CpJ�i��(M�`�Vֲ\ܰ�_B0q�
fk흵X�7b���>(�t���ۭ����"�䉶L���i���W��Ȝ�2(�9x�9.�N���^����"+���>hBN��+>����� }l�6ի�Gg�g�Y@��7�+f�B��Ҕ.�J�|f���!�W�:_�l��j��1�;�%��y���sM�< .M���)2{w�T`d����}%oI\�,�bwz�������[J��ɳ.
o�TAp��t3e|�:eDx�q~Z���ϝBv%xG��{7�2�=@�*B?YC�Z��d�3�\�JL�#�ؙ ��0��b�߂i`�_L�D��̾(��&�����Q�h���kBF{�����|*���0��e��}� �ת�#4���i 재D�ylֺb �X^{tT|)h~A�]�;y+;,�U>Zdt�b��*�ߞ���rO끔����_Ba#n�4-�8��z4/�Zr��E���VT�Mp,����&Θ� ݙ�_=��6D!�(u��z��:�YS��U�_�nW� _%�?���j��s���Q�[)�hvġ��弄��iY"A�a(�k<���5U-r���w��yɌ"�̠��'��t��mx>+�A@��׾�W���qoA=Ҹ'�2|�`1�RVTG��vI^�VF���{���z��h��#�6�+Ġ�� q�"�o���ޛg�d�g"�1n�-qn�Cph
��.�#�DC�9�@H�;Q�*�p`?t���7Z?��)DC5A�ʜ~!�Tñh���\��}�t���0{�}#�PTY`��sbAd.E6r���ރ�[� �JG�$^`�?�����Ö9= b2�N2T�C�m\a!.�;�b.^N���2��{C�<�����#��,aY�:h�=lQ�p�Li��;B��;@r�S`ʸ�R���'%&q��z�N�G/u�%��B����w�}s��%���zG��Ī�s�&���W�XL�YJ�m��a��"yM^� �zo���m$^ն/��m�4�	ʔM@������D��n�U�\�{_�p�x��ew;�T5DX
^ˤ�YȈ��ǡ ����]���(���D݊���G��
����4��j�kͲO������}O��� �&:�y�I8�9'����х'&���E鬻���~��Y@���NZ�Ă{���-I��|���IR�XD����ebPR���qAX��.�S�(��͡n�x{�O�nJ��u'S _��5���A�|���ϧ^)�f�%���ƣ+��m��4�~�9�7A���t���Y�=�]�lG�\�:��z�%�=�H�#�:�K�LOlL]"+����5m�05��(N���L SV!����mGı���T��l�}TZ M��/%��-���;6da��[�@X��d�M���_Ii/z���=��]�3��OQ��h��1�M��!qe�?#�\G�w�Q#J��ҹ(Ms�بӣL��o�ai���i|��9�þ�ćR��&y;ߙH�Ys�O/��Ԩ��v1���%4�m��p�2�Ooc�)�����gp��S�9�Q6f�����N�F��dx�"Z)�*�bܞh&Ѕ5^Ar�����2��lB3S��m��.����2�LOf穎���9�!M�k��P�V���6�v�}����y?���,ΛJX{��$�	(���JrF��#�1���=�1��7�ӛ]�=s�p�q+�/y��_TjI/�4����uWX��y&�`���9[$4/��sk �
�~����J����cR�I��@�^Ĺku'�;����G.p��0-'cR���я� *Ǯ����r�t3�B�PX���Y�k���0}!#¸a�scX>����$��3��op-Y
�t���Is���<��"�׬���/���{�����E3DU�Z��|��Y�D�3!߲y�<�S�,���%%Mx���Gru;.>��0_�%8�S0*Y�b��>�N8P7t
A�+��kA|;Z�`�XRY�Ҧ
�Feg�s"��Jlk��Kw�B����O��isgΐ��girE��h�����f"('}D8v?��}]����g$J��s��+�n�u�ӡK�e���`5���4��������N9�1�h��-���踋$�����6bt4qs�4i������40ץ\�O�w8���M�O���ǵ����y,�o��t�c� �5��U³��~%O��C��\�u1����U9���|\b=�Ğ��bD���Lx�i�M¬ �� D������,@���w9l��ֱv�@uQ���Z�eό�I�W���c������-�)!/rU�2$5�L�l����0�����D�#�����g��$А�Ҭ[׍j���x��e�$�π�@�Q	���� �'ډ���~�� �V�o�.{�ưh-^0AK�8,��>J��hǙZ�u���k-�욁�k�q�xN�s�a@�CPh!���hs~(2�Uo)�	d���p��b��>�C;����l���-6�����0��d����}"�W�r��h0{9
�kw�@q9\�ZR�ﭽޏn�� �ڠ/!>���Y��	+s1c�Sη�p.wGI���ʑ σ�C����䭉�/lsP҇�#2�wbP�[��*B�lW���{ST�@�U��M?���g�5v4r���`_�����\��"�T4��r�6����>d�^n]����Of]Zk>�C��!t���J��xϾ�$���-?YW��j�h�0��� ��շB��z��]J|#D��;��2���n��M�f���W��'�?:��Z$xV��G�¢�Ĩ*͕��U��Wp�]��=�\	�ǩP�}�yWfvɔr�A�U-�2�;bn���t����q��Jqq�k��7e��c��%Aܦ�F_m6�@��)H��;<����ć�<�n�_���1�`��9�=�PC#ޔc��)��"2��Ts$���Ǖ�1��+(�x�u15>�r|Ok��k�ul��9��/���j�6��3,��k׉����`p��������`m�0����j�E�f@6p}��~�?��2d����]�w�j��ʸ�i��HU�����,�rLr2���_Ѓ��"�*�����G5��9���a7�d
Y�5=��s߽��o���tX�u+����Ы	�P�{d��wb��q�Z6��u�G�i���5E�t:$!f���kTv��U�\��Z���9X�T9��!�ΐ�}�} �F)0i�yZ��@6 |lͽ�j��҇����uy�5)T>Ў�]Ux�[�ӂ���ڇ� vc���Oo`@�����5�<Z����=T�D��~��'��G�4�'�~Ǉ9Ъ�0�:w�;��dZ�8-�2g_�վ"��ʾ�Gq�0�V�1�q̋1�'��F;�8��2M������'ic�V�Q�q��/�!i�r�Ҫ��K����(϶��O��O$�#��n�(�b/i(Sh	�َn{�	����h�J�Ww�~;��d�z��66��e3- &�����涊E@e�Ӧ��J�^i�ll����HC�Ĵy�&G����|���5vZl����[O��/�~{�c-�ؑrH?O�~'���6Aԏ�_�sN�a��$���UU�NL.^��/r�\_��󴧖*�54�8/����X�s�P�d��v���Fs�>��L&��Rf�L��~<Z,���%�?��驼X�V���|��΀���FK��ڞ�o�o}׉.�v"��p$\y��j�-�^
�X`�*�?��Xн����x?u�ς��Q:����^�������4��- ���(����)F|2��D������~�_�f�R��3�$¤�
U�U�!:b܀�ӌ�����S��b=4���gߦ�;ify��^��%T2�6�3���}2�o�`����.nn��9C<-��j���|�?� P������%,�o��F�*�	�r�Į
d7�XCs�h;�N<��� f�2=����l�d�B�Y������(�8�=h5>�r����k��pK�Ȏ
��F��@�z�f�*C�L{SQIz��ST���O+�d�<9fi�5�������%��p	J�3�g��yN�!��s��^��<�W7�:�$��f�֘�G-Uc;H�eZ�� ��q"��j�}�%xa�ĝ���
pM�,���h��O��*��纔PJՂ8^\n꠪�����U@�(=�m,�荨P��������\�i\ �BM�JK�{��I�¢��(<?�0��FQm�+C�/�]z���R��On��L�+:�H�ڰR����6@��k�v�>�,i��$4Ŧ��cR�	�o��߉�/�{)G�1�k�O��n*�G�ֳB��J:�P�
������:	g<�ھ�
q�O����E+�-������@.�<������k�|�7�6���}��fi$�!�M	�YF���SǬ�1g�ۖ���P �G�\<"t)��L�?ʄ���~@��˕�q̩�|y���N�m��#��v���UG�*�q����]��:bPU�������>��2Is̙z&��OqZ(�*%���,�P������{��q��id$