��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���~��ZX�NPA�6.������ejSV�d<+O�[,;S�5�x[�$w��Bi��H�pI�.v1%���41�y�%�i��9��伂�i��T��G9���KO|���ǵ�y{��Õ�A�Z�++��e��ZИy�tʍ(��Ӈ�����c|c�D�p�f��d�*-`�E4ڹ�Ҷ���_W��2�PFN����xn4��n������ެ�RAM=�d�1~R�_ !Hz�M[p'M���˂�r�A�X;|J�������
 �y���$38�n��l�(|�Nߜ�P��.����,O(��n�*t��u���sb>W^���EOƷ�/��{j?���6)���g!�>��� S����!��B��������+d�����~�
l��J�4&�󹩡X��)�A^!�vn�x���e97��+�e1�#<���V[�X���@���,{J_�4�\b~�� �XN���U!�^�l�=����QG �8��B�IԹ��ҵt5�p�j[s1�Ό��2V���JSg�64�_l}��S���f�9��S�k">v{���qC�m���#9;���=�/Y����ږ�s��ޤk8f	��1#U�)M�����Q9���(����]u���iW,�mK��+�y��� Y��8�;��,�}�cO��I�G���׫V_������l7�~���ٖfR�3��p����ԒuE=�#��L�����|�Z(�kP\�v�ӓI��B�@����g-*�B,i�����5u�(S�׳�;K�Tܘ\/���Ԯ�-k{��B�"��͑/1"|�0�#�*�����6��$�m�������2�C��]�ɒd�ϫ��~01�H�C#]�M�b�l�{��鈃�)^��
�C��Ÿ��z�xM3흲E[�(в䜰��%��T䨋g���1�uTv�q�o�c�`�8�N�6�)��p^j�D�.TKygxg�f�-��ڕZk�Ȭ� �[VTɴ��k��z�?��͉�^�D������	5' QotnJ#?N��S� �����Y&;r���
;uZ���ĪZ��	PI?-t+�[}EA��Xw�e�j���N�� ���!~���@^RR�<�PyĸC�SkF���d̾���`�)�eЖM>^�r���k�z��~ь�@*�E�g�o�����F�8�k��Tƴ��|��~_���|@km��2ǟ�h�'�����`�6������_�G�Φ*=���6y��T��m�}�k�{K�"�BX(���%���2�?����q/JQ?*��0���sxˈ	�; jI��&*_]���JAN'-�t��X����F�0��6��;\7 �V���B�'E�:�}r_�]�t�,��5���ve�!Kr�����z:*6��K��<Q���P�l֜d���xB=	ǐjl���t��q��Sr}+*�����?�KL�����l�4���%1�#�=�ڴ���tجr��eΝ,+��"�c�?��K4�����F �t| kYH�`�:n�EMjԢm��"�e4�<�b���ȹ��`I�R�����ё������gZ��_���mtk��b��Hw@����O�����V`V�F\�e�`�'�\J8�M� ��FU���+��{���OFz;����hW���V��shlpE�y�@ST�x6�/��������m!k�/*�q�����Q��p�*�� �!A�i�.d�g˨���>+q���j�c�"*�D�b��V��Y����:��%:�	L/R�ph��Ķ^N���,�Zl��刚��D�N�"�`6P��<´�����Jח�j�ͷ*�Za2�����;7/����� �s��u�f� ^� ��O�#�Xo[���`��+t��i:۹�\/�L��!���'/��{���������Ǚ(��-.Y�(��~�Ech�fM��HW�IZ�8����l�J��:��l�?�&�J�ܶ�bg^�t��_(�����`�D!�Ue9{c�mw�TGV�V~�Ĭ6�ݸ��+E�y���1/Wp��E�d��T�
����H�-��NH6��q@j��`���V�:S��̇����H3�75\t�M�)d�9�+�E��#l�0#��� ��`�L�3������\�S�2|F��(A ��ݕ�kk��A>�К=�A��'i�.a���?��-���h>KӺ���O�>W\}�_hge���p5OW�D��{kf�)
oS�������쪈\~����V:ő��;���W�n�l���������I�\�I���\NȐ�����VH���=�f�V�g�]���	m?nbpT��	K_����KL"�+�P~����g�������GNsF����Iq��;�o�&� �\�"k���B��j��t�'�U�A�;3��^�Pf�~tL3Y����ė�x(]�c�P��ŉ�
,O�N'#�v�����j]s���g�j�G0��N����ա׀�R͸M��M�qFS�N��Ř��d���`ޭ-��bd���[����)o�~*�6���
������8.?ȾH
j��{������.���`ms����V�Dc�H�#�I3�E[S��`_G��a�ʤ�f��Zu�wٱ���Z���":���p�H��.�烽�k}���
We�-�N�!�Lݭ�i?#ތ�m��{��R��2!�
	r �G���5#�`�#��[�����y�U�ٖ�b��@mE��'v�i�t�d��b?ԣ˄u*��^�hif�U���!���Y�84�-2ȡ�L������l��5��j)�cS�-���>+���{�Bl6ڕ�D���}X�k��kn���J-�Q$>n�_�g��FR����[*Ѳ�O�J���MI����af��q�ؕv^�+E�kGV�Ɂ��D�x�� $�m� ar+��)��"g�۹KQsRo���d�����.�jD3�⃍�]=X�.�K��CB`��S���I��}��"��ڣwF��\!��Zn�o��H��^����f�=���,}PʨeDB�<J�o��w��R�P��iBt��b���u�f$Fai�)�I�U9t�'���gO�Jp�d�)�l
���h��yA��D��Y����H��)��:#/<���f�t�1G�7X����͓�(bZ�7�9����gR�9N��7�{X�3�I����M�AQ}�	�nqb-.�7rB7-���ȃS�,�MRv�D�-�׬�`߈�q��XY���]%.�N(�Ƽ���݄��CT�/,����ڨ���y��J�_�,(�$T��l�y�YH;�c��ۥ��d������?C� 9��W�t��w�}�H��3X�$�{�����{�%����C��$쟵� ��])�F��w��~�ZtV��*(�Uh�S��9�%���j첔�1U�@�&B1�4�SC�'W��s*��������]s��
���M�{�0�C_aV�-�&�Xr:������+���]�䀮�l����\A@ߪ�<F��r�1h����X��)O��.rػ�y��x|~o�7�vjd�0�@:5C�����Mf�&zSо�c��� %b4U#J�y������zrg���  	���q��O�3Y^�yE���Dm^V�z���[\�2��j9 K�}H��A�ր�����u֔���j�	PhP�D��v<��픃���P�0epT�A7=���ċ�4����C�fnD-h��ը����/r����%EHZ�L�[����>N�<�9m���?�Z'��GG������<.���iE��O��B�*I�ex�YYm'�l��'�뛗���� E��s���n�%�n9�a{o��R��ʮ��x��M�J��.�����膑�rR�L.l���
❻F`s�cK�erj���[~b�Ru���*��hH��[u�B�m.�����w���X(|$-{�b
���y�r�ZH��]n9)@� {�UF���հ����x�ԨW�B+J�k!����b �lGXo�V�/寽^z�Cwp���m^8�"���HX�rn>�wT�8�I٩���nvK�|p`�*�u|�;!������j!c�V]��B@��dѵ�=�*H�X@�h�3�[����}�\-!K�-B邯�����9��Ú��a���;y���.��~��PR��IF1���&I�*y~�7)@��?�E�5įP۵FwGg�׫���	 �0I�gr��uKZ܉�\�a��j�4y~�ҖI$c�mv�C@o����4/�J�,��O�������=#|���;8�_R����oc-Gn��/b��s��¤��눤�1���O�N��!�_�$%�Z��}k�ab��ȝ�,�Z�C�o��^Ռ��x���ɉT"��c�~���9p�̩~V�$q��!��h-,tjfM�[�%Ҝ���	����R�.��`)J���;z^�D܄���+�fߢ����m%&蒡���#�`�2X��+/�b�60*ÿ�0��#���Q)�E.3��/'�lk�������1"���g��x�mi�q���lx�`�L-qR�ᣵ2'��R��o{����n�1�ƕ����^C-�T�w6S!��8s���<حg`�����Ҡ'��At��W�]Е
�]lM�; �>��sT{���A7�@_ז�����I�M)�;� �XX=B�7���)$!oȼjC�g;ƇIۈ���a���3�.���޼�F�&�N��o�jwa���ĲU|��^�T����` ��~��7.�v�����@��(U��l�򺴯��2{c�!qZB\B�f2=�-�Y���V8t���S�"�*.W��&C ⊞{kZO�+�N�S��w�6��^~��9!�_ݮ���|��I O{�f@Z������@����m��k������U�~�lkHI5unܑ'��)M�rX^"��a޵�"�d�7��B,[{?Z�T�b�?��;�1�a�
�`ʆB/��i��7���{K��k�׎�|(��O�����px���`�iLVQ���x���O�u��e�dg^4�"�~+�mB@�4&c �0��D镋>E]r��IJt����mEF5�ۡi��7�,�bn>x�#"�mb����/���ob��3BK�d�6���Ց�����zr ��<�+vi�E��^/�3Y+�?7��pw�y(������$!�M�C��JS���qjp��'G%�,7��їu�cI��)sm���4�~�<��s��m�L��aΟ1��։����dN���'��	�H�x��a��d��Yw��[�(���#�6n_��	%4WL:��M��K����������(&��2M�i�6�%i����[���Ì�+İH��+U|/��Qʘ	o�h��/�t7�$d��ա�����A���XrIX�B9�8�^V����ڣ�:__k����0�����AO�_�|����s�\NkKC�x��l9�4����ʧ�@$��ԍkg�AN�^y�&�����r��g|��+o�._����M����ܦޘ�}�S��H�IJ���YP��Zl�0o��~�����)��Ш���������?jlj%a!�.��qe�f/X�f���O}�H�+Q�-;�p�^[la��}t�&a����I]D���LIF�1�������Oܰ稍Z�h?@;;E��γ����:�!��V��k��d������gZ�4b���:}�3׷?`�\�]hk�A¼�i`�Z��-?W?�u�5��9N���Vr11�k˓�? 8�s�`g]B������j�?�t��0�'TCDx�[��N���`іb��k���#[6.��擼W.�x���:5����,�6�~5��!����ܒ~�k�y�����k��^d.a}b(MŲ���,�#%;6[ۘ!@.%'@��s��G��a�И7�>~�&u��{cfX�o^�¢�7,�u��0��M+cEm67�$�&Z�<ĺ��Oi �Dd!��Cgk�Va�DÕgZye�B��L����������p/�I�?
��E��HPŖᵽ�I��8�X&�����ӭ�f�P�o݊�dy�6�L�S�c/���x�� U�ޛ6C��F�$yG��z�"U
����[�x�?Ҥ���o�E���^\]�|���c�&�������l�V�ed/g��	�*�����J�h�ܜ������lj���Ɋ��/�bB~�s���T4,�wpn�FS�$]��^V��Xe��e5��d�E�|��4U48�n��8gf�������A�-r,;B%�.*N������W�	���d��Y鏮�rc�\J���z�Q��(��΢aD��܏c,;�M����>���אK��ǚ��,lc�͙�|8�C3|BX�����4� ��)=�Y�u2̾�ai4Zgl�|�TWOq��޶�d)`�M8le&�"�2��!v���HE�!و��#�
�����~��v���hP�?C�Ⅱ���ù˛d���Ij4}��@�²C%J�@��0U��~����XP��^����^�:�p��A����gyx��@�JM��2�@c�x3�����o�`�8�88y�<v�m@�%g���V�p>+�� m�#ȱ��cŌ&Ş��7ƣ�x7X��R`K���aD��:�c*��� P���K�R���W��!$�)��[L���I�\��ߤ2 /1�sWy�s[��.�4bd _b���N����ڣ�wTX�z�ܯ��t�9��A�0�ޞN���4t��.�]���jR{���]��v'�'��َF�:N/��Ɗ {�Ǭ���;��J*�E�5Jpt�I!H���r��п�i�R&��[��n��_W´@�
�׀W��]��a�p!2����ID������
��}���uB�u`6�����i(�pq=�"s��ck�}�V=�Z��wb>�x���2D��׍�}�{R����P��
L������0���k�Ȩ�n��D٪L�N��y�
EsٲN�@��5�ef�W�����<*��P��WU�:��F�WJ0]�]��,r]�J��H��&�����P=c�B�Jp��q�~���u&~RTT#�1U%:ø
�'gI��<�U��bv�L^I�@�{�W�>d�%�Ǻ�:����O�ÿb���Ղ�9�g���A�?�zW(�(
}K{?�)Տ��=�T�oC�cc~�sk(j�E��iT3����4Q��Yw��5I6�W<W���Kְăk��f��'l��ߘm�띣{G������{|��M���ѕ� U���a���Pٮ����ʥLDH|�bEpק�Y"��}���r��p�T�t�h� m��-N@8*y�I���/4[�`GpU�H� p�E�1�4�iSQ��S���	�_�GD�ZE�X��r��V�b����ߑn�2]�8rVT+?s�n;����F&U�]ި`v�#z~�	ent=<���L9�� ��"UN��	f�M��ª�1:��NX/���Oys���;���x'��3�_
�}���Q�0o_uyW[��Ռ0�{PL�8�o[����a�r{�� �,�)) sn�_�m�$@O��;#T����m��x)@/�\��A���'��F�}S�nO�Z����x<�n�P��L(H��*q���:�2�OW4lme��<\K@ ��LIҏ=ѳ�������E	�늱����I&.�p�zeJ^*�B�=��}EtԿC�Z������c��d��3ܼ��)d5p���.�\��r����B�<�8r"�N��%�S�����Y5�p]���C���'�NiL��gsɳP/�ټT�R�۞��k] ���.eBC�! ��ҫ��� »���*�1u�"�~��i�u^y��$���z��%Sq^T�����>���������&M��Uî|P'�-��[5��f�J&�Y��<�ad�y[����H��ϧ�>��N�d!��pd��RJ��
w��w/$��%��bA�_�ش�@uo^�U�(]�A^x�K�Q�{��=#������(?̭�<�*N��ư�d��̸Y�?SD�J����M�J�F=��y�7)B޴�3b �:�xׯq�=� yө�T]cU�R<FY�I,��L͌UHw�P�A��2W��6;8C4EE�	;�t��0��*Ha����M�)�a�yM{�]sW�nF���o����0 ֱ��H� j�O1�D��iFrX��겏��*�<��v�˷�N�w$J��T��/$���=����?Ô�>����J�ߚ��gw5$pU̲D<n��7��AD|@;��.z��RS���v��H��]�Kْi��Ő^ѿ຀�.� ���� J�fo�׾�S�S-+�+�WTeo'��k��1
r����� ��?EȖ�a�a������Լ�jX����s���ǋ ۦ.?k�L�L+�cea�K���>,V����t>T	�4�K�Ya��>�����V"S�g��06Uwh���~0��j��AC�����r�� �S���ill�b�wY��Y@�-f_�&*�$ȡ��3�t��Q{�/��6�s�Wf\�Hj|�Z`a�e�����K�|+3��<7�w�}TI�.��a��D�YgrcƠ�ܩ���NX��Ln	n�8�sp���4����_�����7��19)^�D�j����l�ez>�[!\'�u�\s�=AW6mB��s6uy�_=tn�����8�T�)� "��182e4��)]^�ݶK�$��3;c�O�/���Զ.��J<�WӍ���ݴ=x���dj�$��QM�!�;�S��\	�c����9yWI�OH[��Ë=����R&t���M*Ih&����� ���y�F���/W2Hӕ�u�7
�٤!�jd�G�(y���Ǯ٥��$�Q���Ň��f_M9Rߒ ?w���Y%��U�O��k�=s�E�0�).����9sn���д/w1>,̪L���c��&���N.ꘞI�Q|)�������,�N�!�(ŗ��?<#��>߁��s�����1]�
�&��|GC,\�/:��)�:�ycn�D.��(��m�� 6p�d�%Yo{
'��0?�N���$듎jP0�!��M�=�j��{9p�I԰�M�nFm���O&jQP&�mk�,\�9Sז���c�F�)P���k�������'�c�_+���ҫg��]�����OCC�ѿ��S��<�*��	u���VR#Sb�ro���8�:9��HCJ4���^�q��)��%~�P\���~�c�}O�d�	9�h�U�`����tw��iJ�³�e���$Ե�Njt4���&yKq��A/lD�����GNq�G��X}5Ȝ�b��t�'�`���?���� s�=�P�W�';�ɵ�/,a<қa����W_5�/�S��[p�a#���.2YEzL��ɋ��\�S�%�V���i����=�����NV���}�Ta������M�>!HTB+��-��piϛ��y5���R0Z�$���U"�]�p�h|ך�m~�eۙ^����g�M��D_�M����q��EVѥ�D"A�r���;[�{%.>9j�!�VSAbni��P�i�����w��Bc	B�u?M���O����|�"�4g=F�|�?U�7j���.��a��aB�� v�^^�$�acv\T�d��inٙ��Q0k^z�kN���{�@�����u�>o{D���H�i�w� r�f���t��p	{�y�Xݯ$�T�P�ĕǫkM�ax�%��Ջ�Q��͡�nN0n���i�[�D_\H�'� �ku^�e�<z[�w��T�ۆ�c�y�u���
%����G+S��t�j߇x����c]y��Z��r�٘�2eӱE��6�� ��W���AKasX��`B��s�NQ�l��n�4������}d+^�|�!{�j�H^�}py��t�p� ���f����r�ξL�\��D�@��?�0с=&�	����)�����װO�h?��,�|�.�8^a��>�f8��;�}֥�@?�@�gIK��J�_�G��Z+Or�6s\N�����a9��x�}�&>�dB+�Y ����O��U�N�d^�!��̠�$f1[|�4q�V~�!!{��$����X�M5R�\g�-�t���#`�H�WN̾ʗK��ឤ�&�Zi�C�II�W�$��~kSIx 6�$;'�A�Ls��N�s4�bLKmv�]����t�J3Z���0�.]��������<��/��̊���������ܙ��6����׳���*�*޺;oyu�󤚒y�߭�z�����5 r���Z��Q�B��d<��z[+S��<�u��AvTp@P�^�n'L�U�n�<7kTrbm��{\���˾	^T�^*z�Ŷ]�e� [��V����YRc_��\��	���w3��� KI*�|���e�ޣ)m��O���@��]���F�Z��/t,(Cەgfz����6�I4�Mw`[uI]̑�������0�E�/���0�H��4׺Bج>��6�oL^���Xw�!kj<o�1U�֙�#�[I�֕�1���]�:;�/��J��`	0f����ӥ1�x��ZMb��+ӏ����b[��	�2���96ik�� ��������//&�����9� e����ĸ/�3��W$�/�/1��	voē�F�n��~����A�1���!�X�e�Y�*l*������ g� �[4C�NZ�@�B�X���Y�^���N�����t����Wm��&�]0L����5q����l14?M�L=1���E�����&G����[L�����+|�2��xV;�4�`�Ep���q��[��7E? aXW���BP��pu3Q��׽����Q�w[��K\t���G���ݜ4["����u�������r�	n��j�8E�J�
&W������9��&�_ǜi�/���3Ͷ��$����>�����a�[�[F� Km�SKBe�8oE��(�	�-g���T�J^��&���c�ɓ��Ǡ>]δdF&UpM]v!US��M��tr����ݸ�u�	��%�_G&K#"�K&�8�.�Nl�,��ݺu�;�4:���Z�_��e��smCf�<S���\�2]j��A���ar?�H��=��^r,���g���J�8�b���W%��q�B�f��O+.�����?٘Mo����MKF�])���XG��%��nb� 2�I3Bź[e {T���������}w*ty(�Zu����[{U��u�L`ǧzl��{�+�?���Zp�eeH'��M͵R�l��yjWg���S�,����fIg�)��s��F��X�ĝ^2�-ZuN����*��{�d�� *�kx�sP���� �w/����3P�,��<3����+�H&,?4�֌4��H8q�ޮyh`� �$1Qᑈ!tKۣH*������\���8��5��9="+|�Sx��(óf*�� �m3#�\?�;	�OqlF0�I����B��g��1b��,�*��x�w��+���%���W&c��~��ݎj�i�v�:�6R�QٶV汙=��^�6�]`��q�$[��k;Y�*Q��Y�o��Ht9�+�u�BE���/%;�'	��x�`V����������*^e�K�	����q]�h�a��ܲm5�̨|��m���2��X�K�%�I�ݣb���U+�p-p�M�	*%�(|�����լ�덗P��ԍ\�D�&�-����b�����7Ar�bv�!?�R�l��j��^���n�$4e�jl��ȷ�g���t*�B��U���Q��]� 1��1�[WA�4�DY36�W!��)'� �K�*q�\ܪ����Δ b��,Mv.o��pw�����al`����*�@0'8���4# oļ�&,�]H��GW ��Q����5z��Xl�L�E�{蹝-��'���=@.�J�ng�S�3B��]��V>��>�i=����F��24(8}�(e�;�!�vlfAp�9B��2����P���B�a�1��F��!���b2�����ҹ���5�`�A
v����v�� ���*O�钠s.Y�	i�Q	�:b�W_6m"$��MjTSg_�3sZܳ�����A<&2�X	b�bR�?h([�7�Ź$�@�`C_���Ru���tzb۳@�X9ص<���<`�`Ҡ��F�����
B�~�~^*�v�t�@ɘ�0�/`�0��y	�9ech4��t��xV�f��B�x��n���!�?�b�>b�|��B�wc$���摨pO���?����(ڷ��Tw�9�~���)�\Wx�X�c��?=Z,�������@���/�.j&��ߍ�0��z��"���H�IT�_��E0Shn���A���H���kr����CX:b*%�,���b*�\m��FB͡��B��%_����Cg�	�	evƎ��b�b��5i��z;Z�(���QA�텈Mǘ���%G��}Bە�	�����$�>A�(�	���1��|�o���߫�~�6��D��]�h<�/�V��Wخ#���;��H��.����g�XC���*�^��s�Ҝ(���K�S˓ï��7)wu�+#� �����}n�V��P4�W2��`B����"{t�x��7�����R�6�V�6��1`���m�_�la� !U��4�©�w�]M��*�B�`^ ��x�����<}Q���]���V��n��K�	H)�9�i�A�.z��qj��o���a��0�d��]k�������g������j��`�R��ܣC���G�/HN !Q伔��^G�=�{�'=�U��rձ$�K^��U�p��.�\h���u�����*F��̵��ɡ�ر�t��*1�)�v�����A &d�C�a��ޯg�9G��F���G[�߿a?9d�pѕ��W�%hA���1Wq}����0؅9�q��HW��=v\�3Ds縆> ���� �0F@����V�܂\��k�frW���B�I��{��2�1���]sO������?>�%����ĥ^T�~P�j��wÑfD�����4S�*��@�N��'�mN�sL�Z��/c�j�Y&�z�L{����.muf&���g���y��H��-�W����L �����.�huٲ��%\ �73KZ%�; ܢ���BP~i;�hv����ܒ��H=��>p^���͜s\{�o��S�R�}�4Ug�\6�:��?Q\�]��L{W�|$�/{%�R9�QVt�Ã�n>x��!��J��S^��l�v?a��t�0���F���|`x�c�����*���H���*����?���x)l>0[R����qWL]�DS��X����g�Wb���D�=�0���_��[�0�|�\Z�<1d��\���D��7�����ߤ���j:�/���n�E�a"���
���|j�N��dK��;��q��.~}��]��NY$0��AK�m=�6�/��<�c��Z��>`�F(��Kn�A���J~��VB<�qZ`��@��tUr��w���?;���M��ۧ�ur�PD��,7/nh�ͥ�b	�Veȏ�*g�X�]�I(UBp��I�,5���I\�>Y�(;�{%w�!1��_��Ź��c��cR��<?���-g(��e��O��g.+��R2��Q�*�]pߴٻ�!��_�Md��t��E��,΁� �������U|^������&�&%�r�<7S@0��P�+�n�d�� ����Si���ͮt0�*)�i��M � s��Pt5)"�	C�f1�WVM�R�T��%-4ǣFܲY6�}A܋T�
r)~(}F����4������l�-U�O}��"O:}��n�:_oN��U������yϰ�G8��0���#�*���*>��)ĤR��B��Z�r��5��	y�҄����LZ��M��,*�@-�*�]|���q�H�d(� r���Yͧ<37��zY�R��Q~��9����,D�/&غ�����Ѫ�Kjj�5�a�)��5�[�TJsOdLK������#�M�$kI�5�ǵ����5���v������"	��䮚ÑNA��]�����66pqY�&2�L�$�k�9�G���7�;��5�U�YN���L�/��d�9�$�v� �h���+����c���:@{˜J��4y�=<��}���ळ�6�8^�qR%W��[#w��Y�~���آ�-�7����Z�O�����n(�tU����k~��yB"�f�K��"��&��c`�LT�z�UpHpF���%��qd��e�sa�!HH�}�\2N��~1�z�lq�F�g~�#�x%x���@���qT�NQ^�(IϞ�CM!g+�a�����ᠸ�������;�Tw��>��Y}q�S���Hۅw�H�t�P$!<pmA'�:����0p������&���Ƈ �6��!�ލ>�T|Ee�3�@��X�s]ɑm��<��}���%~ �����~���Dؑӗ���ilԣ)^OHS"���Ҝ�*��m�se,�6��Rp��%��<]�u���t���]�����Yixn��~��`��'h�B)��Y�g|����?�����r���ށtH���:`Cacg�6�3���`Mۑ��˵��2N�X�%���1�U���;.��2�#!f�EQS�1X�)t�)�qIzA���%��Q��IΖ�/��..I���b7� ����9*8�+_:$/�$F��>&��,�3�{Ҋ���/K�Be���
�i723�����'c�
k��a˪`���<����R4A ([���aM�TiC����;�e��g��B�r��D��1�L��� �/p�@��M��~ff6b�6�)����������RQ���7ˉU��H����$<k�D��j�K� ��d�AA��l��p�ϥ�c�hDSF7������I#t�I�-c��;���Gd���H�LX/ۇUL�x�[�mK�z(��tk� ��4Hf����	���z4V�N�=M��h-L㋫W�N�WL��NM��9�(��U�����y3�0[#gŇ'q�$����b�]r����x\MQS�j*Z��ɗ�쉰+g�S���>���H����o5�J��vr�.�n��c��K�P�MNG��]��{��;� ez:�߯o�X�����>��r&�0��R���B#���5��ți)Tz2{��� SW�d����sWHbY�y@����xƖ)��g�A�����
�yi��E���6�Z�����C�{*�y��F��?��R#T��Hm �u��� ��)S��u_�g��տ�!��@�on�1�R`����4@v0�c��2m-��������&��م�O��;"��bĕ�X,i�"����
\��?|A6P&�i����/~T�BYa^L�y�qU�Ҏ?թŴ�x����{�d�.M9�����Bc�rCz��	��ep���\n�%��D����Ӣai�A��thmf ��2��%�'_"��<�
 �˨a`uR]����Ø��5���ıN�mU; ��)���[�V�Z1c\��1*����(�|:�C�0y.|�b�`�0�_a�)H7`F�(�^����a��.P�e�>"��*әB1�L	3QGI�����:l�)�[>��vR�6����G���������{�����ݾLiX#f���yl�F�A�]n_����{t�1�s�}��X;�Y�/�D�p�lT7ZF��b�Я
�c�Bſ���fDL�g����V�_V����Nlp T�ߒ��I�&�8E�Y��JI����1�-Z�<�5�Ŵ/lB��p	D��KFW��N���;��Q3�񽡉����9�)N���ԻƂ_���$����k>�� ���g���a���x3�=Ia@2�ں�*��O��P4�:����r�	6�G�'�w���ԫ��J,D}�P� \��û=�u�.uh�/o��+��؅�?r�1�����-P��&X�>Dh��kt�C����]擏�@O�<,�W�^S�g����d|T'K<��~�K�jٜS�AG�����_��w�|��"ܬ���&+��*v�l�����k*���^;*����]�s�&�,R�̙3\~J߮|ui-��6��)�7���$6(b�M����g{߼J�r�w�$45�<��W������f!�BeP��doJ&��[X�@w��xݨ]�(8䲙e�B�=���;;��1��[��7��J�����K�Q���B�;�[栺Tעq:JG�����OSؕ2�`����X[��m��)��￵�Ֆ�κ�4�ɾO{�������^Ag���KLw��^������|ǵ�}}�yv�e<�0�� |�}2�P�=dwK!)τ\ͩV]���ngdM�����6_:�9ߥg�t��?���&U�xv�C��J-2-H�(F3��8��H�Y�����#8�<^A�4�ڱG��+��ʭ\��-pi����T�Y2?�=ʒ�Z�hz�0L`eK����&�U���Z�n$�J(po��Ě��