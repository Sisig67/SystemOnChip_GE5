��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%��eW�z`�.�ThdJ���
s�sȹU��찐�S� ���{$a��[��ѝ6�p�>G�\�א��,�:�ڪ��.����_��/þ	��{�$�<�jY�_X��4'�]��/�(�5���Vf=���)���tǐ�G���ag�gL�PƱ�]`SY.Ȟ@�2����e:��_��8P�LOj�l��#j=�F9�5�|���Iz����T��ӭ�SR��.6 s؈q�j5[l,n���K�6l�����EF�/j.��_49�MS=�A��Ρy_/7*��:�� Y�Ź����W�_�&ȼ��xma�+�0ov��&�8	"�O�Ǧ��j��U�|�rF�<�e�J���K.%4T����� q�@�Хݮ�TJs%��L��?Z �^�-���V�Nk�\�{������Qaeܰ��y�(_��2��Uz�0�Ō� m4��m�)�wD�ٖ��o��gԹ�M��ڎQm�G�W�8h�U|������<\gm�M=�@T��oY��%�� �ͳG��	���>�������w
�+m0\�f2arp�A8��_�~��"�0-d�Aw������F��i���(�F�ճ��| ������8fT@�I\��D�R�ڄ��,b��#/�YAn���1��y��-�q�G�����'�QwYz��x�6��A@�q/��3�;�O<�U?�˚��6a{ڭ� f�/�d�J*�3�J�w8@�|j+��^�cB��s?5����4졁���N�(_͚���.�"�[��"m�U��״����5�ʦ%�%�n
�ˁ냒�D�!H�I����.Q�۩�~���)F�y-�&���*�No�i��������l۶��BX�G�fH���<!�e���(�%�mPtĤ|��L�����r��56g\f *"����ű�/'����vU �nPْ��p�\����'����栛��5>CW%��<�{�3h���)���P��ObD�!���(��{t��Ɗ���m�)�?�݋ą�gtv��q�*Z������_wW,i`��*Z��^3s��2z�I�q�jnk�˦�~6w�roa�Bɖlt��
��NR���"�2�~���@3�'��bhU[��TKB  �w�9��L�>���n�	�g�y��Ԡ�қ�Q�w������K�����0;r²��K�L7�w衚x`�c,��@��� ���#�&�*�~����D��vS��<��㩱e���nA� -�(�p��˶����rwT?�5C�W����_d����Q��E�y����q|h'�wz;�O�rm
��3M�!G*=�#\��h���i�'�@W���<�1pW��zGCRb���e�u3Qo;�]���(����N�Ͱ^YzڍM���J.ѱ�1�����.�v��l�>B���KU��I&゠e���\WX\!��M筑6��şȐ+�jS=��~�%ͅpy��<9�*pNHn=fr��I���v`�rx�N�Q��g� �Ƀ4�.D0F��rx䔂�L���������}nJ2�Ʋ���H����s���֬����UØo|�����-�O��b�D���%B�`(Υ��B��B���lIVuĲ�ą�5�G|���X��T��]y8��]m����tV*d:�
�IY�{�[�4���kE��~����K�E!Ȗ�xC�
c����F�1󺛻ĽOH�4�G�J)+�L��/6�gl�N�f�����&kY��ٶr�+���zUW�Y(g&|�W\� Q1�&�J���&t*��]��=�5��r�4A18�Mk&�喗eƪ��C�����
g�\R�Jѩ��RǤ���
��+��r�X�{�pҍ�>�zY� �0����s#K^�� �Q����S���39%�l�{ZYd����o(��ғ"2!a��ol5 �&�rw��W<����P��޸�»�Y��"v���ɶ�I`�P�Z��i��[���s�b��
�	�л�Zbm�:h��"��M���?Y۴7�F�[C��Hy=-��+#�]%L�����$��w�����@�;.yu�tɑG���?h�^��1���ˇh�b��s��i��7��ȴA���-��K��5�ύ�Yd׌�{@Q��'NkM�DN�)�������B�@�����a����ļ���	z�s���C|0$�?|k�G��ͺ�40!JNl�IM��6���q��3���1�G@~��ζhZ��V���卻}\�,����r�e��p �;��0�d�������:`�աv��F�k���}f ��Ei2�-ƞ�O,!�"k:�Mٙ.�K.q�{`p�[�}��l�d��W�hE��cvu*@n�I��}XK>;%=#�jh�A˘`��Ů�����s,���q�?̃Kf57�1,)��,���!-oO\���~c� ���A)��p�]ɠ��){��8��6���w��J�����[��Ui)�i*΃��
@�ςN����7sbW��r�x}�7� /�?_o�ā�TklsZ0�˹ѳʃ�-jh��:�i.YP/��kQ,K8��H�B��b������DD��X脃�vȦh�<-�?�T��թ��HP0�S�XLЙ�Y��=r��gS�����R�-��ƋH|��W�T��9�!dќ^�	GA׸2s+�5s\�]h+�6*��y����D��z�r7�8Q�q�L3�|���J�\:Cz��^X6rFʄ�Q$v��.zi�oj�6��������a)6"Up4J�fwT��(n��Z�˟��Z��N�����/ku����+q3����Q����*�֤�w:{��XH�B`�ڡ�eF\cRl3��,PZPI�.�$����o+^��`�p�";�D���I�-�,j>o!3�ߝ��wJ��7|d�6� F�¿�����CF�D$8|�	)ȉ�6CȋW�eap S�#kh�#H#�B@A�.pW�nc-m��Dw�5ni�D>�9�7�CT+X����v���}6s��0:�,ᯩ=yS�%���C��kM�@?A>�/�(��g0]܆��5ݸ "�L��g����L��RJ��$X��#����.���ن��l��C ��+���N���X��qn^�����H
�׃����IIC���{��h�4�{5M��a�m3�J��� e��$|�,o9�;�޹?��Hu�U����|�����k=R�~�>��}<�,|(�R��$9l����ݬ���*dBB�b���;�_n�oA=@ͷ���V�@,��������m~2d8"�<F#.��l����4(}S����.�tw�bX!��ߊg�y��Ϯ<<"!򮞦�S�d%�J(RĚ���u�9�oN�f�����< �q��o٪��O��?���Ճ���A5�85��4�::R�yF!�6��0� ��%F6-��'��v�ٍ�B��ِV���$4��ki��qBvZ�p+�UsJt�[�[�#��
��Zq�FH�HF������+f߈(��Le$���q��k ��ݩUL��?	�[ɀ��`=��n:u�yd��ˮ6�3"/"e�&�0��o|�o�JV�1�Fm���U�� 5���X���&4�7Yg��� M�Y?��$ICBdH�!��NA�Fuu� 5�RLZ��)mRj��J�.�x|��s��a�߭(U�zM�c�S��\�� 4��C��"v�O��u�Q2"���fB�T�<���"�/TA �ľ��M�(Z�l)��<;���o]��è��ԃH��%_��v�u$ o��5l�F\s�c�����f׼��J�!r�~Ņm�� -EF��}d��Xb�"�l��q�=eD+��=���4X�H�r�~��E������7��r�V�$��L�Ξ�Z]�F�N���Xm|�_O"qޫ���KA0<ˡu:���y���)f��V���������ӆ>Pz�m���pS*Ƨ�9ijF��33xe�.E�o��̳|�c�ܾs�=���J��9�v�KL�\����0e�e�p^Q14[�n꠹|>� �1�$S��v<C�R����,0�U��k	���������$�ިC�H������줭�[�qi�*`�6 �������W���vſa���@r��X�p��=�%����b)�Y��g[J�	:}�]� 7iM��4�Y��^+�L���r�)c���"�e�<�~��6�J�y
�\rH�4o k$D���7�_ �?hY���'L/�u ��M_/��1���[jV���>���Nk(�[�e����i
������l�$ ����?<��*UG_�&�
�δ�6m66�� �q #_u�'k��o]!� �����'+�Ld��K34��8�ʴ�Q+>���/>��
�9}U�np%�,s�!����U}�;�+]�AW�/���gP�E+�\X ���]I�G�'�/�su�#O�FFEП�eA���i9W�>��x����8GT"�l<�d�L�����3x��9Iz#g1�Q��i�Uhܻ�-q*�i�
}�\�XO��&tw��3X�����jl�yk��S��T�/E,�J�d	�1�mwk�^c�_�gc�R4}�C|m�� }���t�C�B��q\)�&�a柍�Ⱥx��c�D���^��<h�_=J/�ti<]�.iZo���mA���b���c���+�C�ٌ��_��
S�����n��5��=˙��iq�cK_�"�`�u��brPh������U��l�Н]z1����}��ߑ�f�+:߈ݏk��3m�W���h�ۦ`!��s�Z��C=K�M�
f��wå�ɦ���\��V �ߛ�%�)��^��c��?P2;"�Q3�O���z�+!���J�p�<��Z<�Uξ��S%J��9��fS"Q�Vv�����x���w�ہ�|	dz�7j�=i�� n{V�G�	R0,"u+o����n�PrTT^�ʐqm=S'���auߴS,��֎=�5;3Đ�u뎽�;t�KGi�i���h� �=yyY+��iH6���=��15���2b���/8��IHyM���m�J�B�*�\���,��j�w���`�wj�{�!k<9v��7�Ljuo�u��l�I�H�j�f�Q���h[��I���?h-��~_֜
�9N�E^)���i����� }U��u���Ny�_�^\��c_�+��b�r&�.V�AR�C�U��n_��Ap'8���ݎh���m�K����c�dr�oilM���1������("�].,e���"�`��� �͢[��턤�R�zNP�΁�e� �8{�mq�3FZ_� w`)3y��|��y��֛�ί-'Y�>N���M/z���i�|�>fJ�������b*��eǿ�P�\̨f�'�/,6`�7b'���I�7�eX(>�~Wi
	�%:
��[�.���ւy9vǔz`���Ia����9*O�+�ؚ�D�W:%-h�ˤ
룛x�2!��/����!��� c;M�XM�殡u���[�* ��g� Nȁ��0*ϛN|q2�i� ���>i���ʧ�
�a��,�r�2�c�!͋�	0G��	!VXL���V]�f ��<K/��qV��L:�u��a��,�W���$�������>��U��RS�@|��[C0d����.�����6�[M�a�b�=@�@�pa��W�����*�8�c�9GZw?�Q���n<�`���۝>�A_wΌ��80N�=��Goyx�U�l���m�����$u�1����[�H�v	�u�k��<F���*S��4#'6$���e%�ܢ ˀ0�k*Q��M>�j�M�})Q��h���̒�K�)��$G�Ђw�v��T�b�-��s32�.����l�S�b�o�з�ۮ�L}k��}q�,�}�����.v 5I+'�+eЋ���(������},׮�6E�Z���O%ѧ��&����`��a���?��V�t��)qK{?��O�� �N�u�@���y�%�����&nK��H!6�`��Nc���v\@�?�������T�-`q��M�P�Y�f%���t�����W����b��Vz��ux���z4�P.80����g�T6dS��1.ʈ��?7�q$��X���e9��Q'�t/�����2P���uFT�C۸}���N�{c�ܹj.�����k��s7�?��u�^'a�7e	<�d�I�#��4ނ�rU>t�MM� r���z�8�Χѧ��X��+T0/�j�3�1E�:�h'C�$Ye_�m�/���T�j<Z+�X��q~8��ag���Y��A�)h�	8r��\��0Q?Lڨ����7�$���E��k� VuS�<��{_�%��D��� ���A��t���4�Fu���U43�_�ʰM��tYIF��M�W��Zu,6���sU����Ԉ��D����w_��7~�xY7s��r yt�W#z�lᩒ1w�ךl4���4�XT2΅���،`��Y\�S�����)\��ᒚɒ�r���"#O��d��b?�Z�8����m�K|���I�NƵ3�؏��i
C���K�<�'1A�w�g�d{?��2������6(��xE_�P��4�������ό�H�8�ǌ��=a�ָ/:���� ������yxpLLU3u/���IsA*�֙0.��I�a��ه]���,@/?*���g���X�\��S�|-i�{��$c%���槑.�'|����0mǷ°�H6���|�D[\g�A`y`�Mu.�^<|Y�'(&�EE6�9zvur��͎�t�E�:G�Z�I�VU |�˴��H"k�݊I|۽�{�1�rF�Dx.G��%���*�W��^cXŉ��C&�z��6!g��q�+"�I�]#T�`8�������+��,�l�
�\e���૪����y�II�91v�a�N9�Ъ5�����4�Z�.{H�x����3�M����eY�?�iÆ�������U,�۱��C�o��,E�m��ȭ�E��#�.#�)�����WMs�蹷r�1�%�qց��L���� P�"��T@�!	:"�C�;�<7�?��������`~*�+�������"�BK�R3^/u����֒Z���I�c�l<���+x�۬=vA�$y�{��(��H��'���g���/��k��N �ݣ����dDl,I�k����^T�RX6�P���c����67�S:���R�%�DҔ`���hF&�!ߢ%e�G�Ā��V[�غ-�Z�I�6�;y���-��?���Mz��~˃]U�d'�s�����2K�?��`�[u�ϸ��#�¨����A�$ɈnVW��RQݲr�x��?�ճx����Yɳ���P"�$�w�Ԣ��G��%R�&2��$s�+V}s�3���+��g܇f�3n�wըm���/Ǉμ߅�ôVl��_�ye�1�YR䝎�+�������a�y���J��*U�v�N!�D;�IP7���b %XUY���/��=Υ��Kѳ
���C��.���yy�oѡJS�bbADRb�ل�

Cc� ���C��S����q� =J��澼>'r����do-L�W��]�N`�"��/�q������-9��i����5lu����c���T�;���&�ݷ���3]������q���pߍ�a��bv�NI��p��?Ⱅ"����@rh�ċ���\KX�s6O����-���)��9�ϫ�aQ���GK�	2lzLd�I������<@`�h����r���Nc�I��D�������2�����H�������N���/`lmΟ-�8����{wf��R_�0P�[U�`�liñ���y7q�@Gl����P@��q(3D�`�����_}���Q�*T��a����+��()O��>�# �����6Y/Z?E�c$#2�@�`7DD`2w�1Q뒎�(�����^�<����[�vv�h�c��@S��S�!wN�r�\	�do�4����#�bp� ��N��J��CB�9�C��Ur�6�dp�K/	�`�eg�O�>����pî`��bh겍���:T����_%�A�?�V��Y�yD�N��R�o\�bSC&��O��9³���!u6�ߎ�9���L��gu�_;b�x'��������UQ�li�<7Հ$
�����7��g(�0���3AՋ�&y_�3fO.�.�e���X)��ĥO���<���Z+���C�����X1��+�7��GQ���d�?t�!1���>��ݢ��Њ��O���V����K�B��N�MS��~�LtΧH��S���!r���kH-l�X�G�/�G,}W��F�� �=�w"s�Z�c�k��u�A���0۽b���;�E�|>�����}&����<��~�K~m����'	SZe���#*����=~�T:Y	S��eϥ��V������Hr]�i�7*�*�z�(�P�r�,z�\3��RIN���&�%�z�V
et�ԫ��m[mxfHN�޹�ۥ����W�Vs���ӣ�J}A6#��&C��=�=��o���o�vP�X������3!�w��V�;;�����U��Y�b��fO��ŁP�ڎ���f�����#X�����r��׋�*�g�lQZ;�X��v\�m]f>E�� ��]��y5��g���M�A	>'g�M�'�E!w�H؛l��h�Fb��3��̃�҂��<J�H-���p�v���*[un��$�y�&T�p~������+SF2�E*����ٯ�������������qa0>��7P��l/���,N���bԿ+��j��2� �qƧ�;KH!�QSh`I\�����^�j�0�Wq����7��oΆluK��aF��9lu���f��������!�Z6@#�w�k����Ȉ8h^�{�|�H#�\ʿ�ɼ�BS������~�6��rȏ��8�ٰ� |J�����}w������7���|���l>@��l�b>�/_�]-�"&�Gָ�o%G��Ni����>oKc����p`eW>�MN������ե�2��e�GY�
�R�p�["�&��5�Ռ�0
E���#56,QW?͵�	��;��.%w_��}X����ܳ�EN�Oɡ|��5 �SW���ل�m�Ș&6�6�^����ѠA�K���g %�����2_1���D�5O�"3�ܮQCA�4e���3,�[n���-5��U�����}���W�V�;���'�$m�:}�
��>	���~������>6�\W�PW�"���PN��ځ�n��Z�4�N̘{�F��h�O�^��B�FJi2���	�@�M��mЪΓ�7CM����mS'�|Xx�?�Ď��Թ����)��(�8?�wlT����F�Kw�s<�����
�`�%�G m�XD���h7n6��&���7� c?fs<�?x*���F����(���Է��p!����qjD�wE���ͤp�B;��O����Q�!!��#װH3�����>8��۹�I.fh�m_6P�(�:x��v~-�[�%�5̻�]Ü�v:���E��a���!	E�Kz�d����z�������^�W3ۦz�j99;� ��`e%�2��?hɉ����֊��1�f1KZ���)�QK�$n�oR\�m��Õ���.��1����Wb�o���A3������*W�/�d,F�O8l���͚���Z�k2����!�V~q`(�0��w�ZuPdl]��fSs��W�h�������r�����
�i��ǩ���'J}k�*s����[�wDR���l��=J=�F�ѕ��wxBas��]����x
	�ٰG-6p]}V��~��s��L?Ͳ� m��f�9ژ������[uM	�s�f�EG�m��"�e��]�����xa4}`�����K͡�;�Xح{tMQ��M�S*��c��V�i���ݢ�D�>���:B�%�V�Y=�H���֘ �B�n�γ捩~b2�@쒘iZ�Kcg��n�gO�pf����ȩ��:�V��	)Q�{u)���y9{�ր��Ɏ��B>��h��_vhx^���p2W�Z��OdZ9�xq�lmG���k�H�a{������>U�dDye�u��;�TL�d1m �Ej.�ћ����o��,Ö�-IP�hvfw�p����0tԥ5�5�^;�CP���`×G�'��mH�B'"�/Z������3�3�,T�]�w5�v?׊X�6ˀ��F�MV��sv��8�h�~�0f�h��%G��X�~���S.�^��6c����lx���V���?�n���1��Y/.Д�>4�/qY�BAP /"��5¸8��^j��Ѳ��g�Խ{�e�I6|�r��on@W�l��O:��ѐ�}�I�J���g��o�Kȉ"ҏ� ^7;)תh�9tW��/j�!��[G�Y�l������#.��f�}UD8�����x�qFa:w��3^L�o��m�=��b�
�>����}:vpdS�vo�N��W �yM�,lv�3v=���H��}lM��/�O����$��ܐ��Nl+ |����z9[�&�1���BXY'�؅��7�Q�Q14z��S��/�h��x�t�@H	鑡T��}��s���~?�������K��0kw}C��ܲ�K���WN2F��H"�@4�My����gd�C����ŋ�ruڀ�"��ңy&��@���׻T~���^ �ڂ��h@#�]q���=`h.��E�qA��A.�$�q�WY_H�q��<S�i�q�yJ�V���`3�%�Pu��рwd�>e\�������w���qk=��^������߈j��u*�	�M�������S�gG��^�=�&��Ku[�z���H]�h��X�g
�L/��g1%"�3O�;��l7%��a���)�P�k?����=*Mɀü�*A��.Mv�ړ�oH�!j�\�Ʒ[{2Zuz���ڣR����a�Q��_l�)�]�t��ވ���k�L+���y6JU�L���6V�0����0���{wكץ��AK�;KP�ga�Mi�(�`0�-A��v���9���c���Q�V��	Ó���CĊ~]3�mQ.5�W���1DA��㍼�dz�mȆ��ڏTVC�_y�%[������;���$�T҂)pC[٥w��^�v��u�M,��p�[0Ų�"WR����ߝp@9_F1��Bk�06W��E(B�y�O���E��}<�#�Ż&ǏȎ#���Ҋɠ>r(<\zW�c��9+@�x�:��N@7�/��+��RƦ���KF�΋�5��X�l63��1/J\���:;�&qxW}Q?kH|�P�ճ� �G����il���{٢���[����IK�� n�?�?v�^������Dc�}�����h���Į�����A_M���ӦX���=!W� U�h��b����T~aA�Y���3�;����e�})��AO��^[�n�RQeL;��7Q��s�:����� �.�5���>*'2̒BR�8՞u�-
U�c��ᅈC�z#��{GP�1`�DW���>3\��na���S�P����gg�2���I6�W�d�[���^�rQ��،�������U�Xߣ{lC�X-M�ܤ �9Ν$����/��Xi��#r3~z�GAϐ�s ��Ԙ'����IՓ{4�HH��6� c���s�������*���B9bMf8B�ӁX�Վ|M�ظ��K���L��DK�E�ɤ;(��Ѐ|lH���	k	\��B)���ߙ��R(GG(�&���:���WWD���VX)�HDyҼ�L�;/�Ą!�C�	QVe��s��`��o'����ha�h�G�Z�a�1�cI��)!7��z4�����Mg���L5|Ł!��C����ȱ[�g�
Zcl@��C-d{��Ammy��զ���r��r*�p����R+nܕ�UU�r��K�;�{ci��-b2��!69���w  ��kαw����:c�6n��jt���L�&se��l������~2}�{\?���К�9�!G�����[��˺�C������͔q������q����Þ���Y-��^A�	L)v�D�uBT���QJMu�����GW�B5tq����f.W��h�ݨe,��̴Up��H;��;��{���j�Ŗ;�f�SwKt��6��	:L\���p��a�L�o��x�V�Lqa<Ϊkp$�h�t�W��U��*��{�N�;��$�T*�i�":�q��QQ��nn�Q�d��9*��FWr�?*r��&o�f|����~v�var
}�t+���x�v�,�H��o�&!�h_4�"���5f1F3�?�9l/n-U�:���8?�Z�5�G�k�|�_��V���Sl
�|w_�aJjNrs#����I�"�V�پ����u��\\).��=%�`%�f� ᨰ�)l�*T�G�%M,�K3�Qa���S`k�*	?_hAf[+���~9�,*�����{A�9ԫ�D�+�L��
��t���}	>fAIc����.{����w���3/�9���9RS:k�:d2;%W�"{>�#G��{��u�4����2i��5��b���ھ�)P����B̯�CJ�Xq�~�-w��96�/�y�ZS]㢭���w]�W:�c�؍Ñ�^���x����8Q��1�,��*}u_��Y�F��ܺ����j`ɹN���r�^�m}fH>�H�lΨ��"遮�6jP�Q���Uد6�nL�J���a2ȶ ���a���)�p`7���B��w�n6z��!�j�dލ�	������xo���L�au�=�w=�QɳF��w&&��f�/�*`�4�y�P�Αfy�#_E�5�����+JN�(�ֺj	hNE�6��YCʽVs/����TM��N6��H���p�%iΥ�Z�v$���<���.��@��¿�f��]|�?��S��]]lg���t��7���������^�k)�3K��6]���Z�#�0@��,T����//��0��l�������-2o!Ǐّ���?2���g��*�[Օ2߁𿞓ա-�b�牬���!H6��%T5��8�xR�c�[5�iuň`�><�F��s��ɍin�z#:�(�q؁sz��N��$F��[�U$&�{��t���;�HR�A<��J��X�B�]&�~~ 8�Gd�RE,�����уCy#�U��u0G��!Z(O�$�#���M�}Et	"0��N��`02 ߻�K���N��h{8ebI	�񑻠�F?�Ψx�{�p���I�������������
 ����r��ʍ/�w
)�K����.�������b�����w�L�銧az�B!a��U?Gw��	�p{��h���<~Q ���ݺ��76y�u���.F�����t%��L���g$�y������1ﾐza5��d.�h���c5j /��{�.�쌏�ŉui�R��W����Q�^jbc��ii�&�"�L��1R|G��T���D���d<�%���h*��H�λ���������I�<�vY"�١�.�k�o��:��*��%#��/���UY��8,�k�}���5p|��{Z�%�7W�	�t�݊�L�W�S����_v�u�F0����b�������2%���KƎ��n��ྋ@=#�D4��P�ZԵh+�._*"�C|�uƽ*�'���5���������n�Y��C��������#�4�J<��P��$���V
?��i/�gݩ��]�35O�'�a�t�����<h\�l��F�/HY9��xhMw'Uu�MO�[�R��ZY琍ʦ����v�=>�����i��{U&z�4���h�m��i��[���v�(6w�n	&��&I�'\��d�]Q�h�RE30nU--i�حMC�3W}�\����?�����s,�v�� �"c�I��ۊIg��@$܊���~�3l���>��s�&�1Bzt�u�~�B.�]�Ƴ�%�^o�	7Os�	��K1���6_��M͈!�N�e�M�v$��2P!�j��Dr5��x�ƳΨ��짷|���Q��e^�J�x�P�����g=ߡ�/�24�HEE�U8XP]|�S�m� �5Ӿ4V�������գt�߃i6M��/��g�?��!�E��E��T��!9=d'N���0Z�����Y\7�|iZ(/�Hd�B@��1�uQ�%�����#�$�{�2��-�kw8�_�y�d��B�݊���V=��oUi�ps8�o��5�� H�dl���Y���yz��O~G��H�ޱ��my��4�PU�����U�h��@�.}�iy��q?my���͚A���Ŭ�"+6�h6�� ����4�{	���g��mY&�&��;V/,���U�V�I���WQ��.��F�
Q��*�Q�	���{(���F̡vͭ����(Z�j2u�kߐE8�:�s���4�PR�v�E:E=�B�4��y�ꮑ�e��iv���ƒ˃����A��,��g_V���x���������VYMC���}�ª�s�Paįc�-	�Ѵ�҉�,Q�����Ku�^0��>�^l�+,� �����W(��=��F�ń���0���?�����|� 35�s,W��j�d��p���;Vt�f��U�i��9}��A�SB�)#Ml	���9������*B�JT�Ꭿ��r%���
v�U�i�1<n������9��|&�H�'3ֿ�HU��;��gU�����H�'���u.�����8	�<����4<glz'����q�aJ�s��Xi�7�L�%�+�D/�j_oVfhB�j�g�p��s�~�/�K*R�I2`P6���I)�{���E��g�����X���d�5��̬+�sLܰ�:�7��pa_\���l�/�?"*O��%��j�"�����f@�ӫE���+���� ;��������+����$7袠��x
��;}����m"�w{��ˑ�` ��O���H������Cgr�	V�| 78�"T~��|��Ғ�8g���0ȚC}zy�'��f��ؠ��.�
	_�y�y�צ�ij�3�3�!��k��nB�r���Q5h����mv�������[�|�����U�𒌢~oy�'e^��-)L%mE��=ȱ3k�F[1"�Y���՚���%��@�D&��m�j��HW=iO��xr�+WE6ʶ�Q�E�e�;�ҡ߿�ƃ�حJ��}ԠS��I�O�7^�X
3OoS�Dx%kf��>:���O˹|�SU���;��{&�ܬ���[������t�[��ϭ�v��o��Jo'(�9���΀�������d�������a�~�/��
D��\�^�#
-w>���;I@r�rF�:�l$'�a}��>�t�*@���`mh�������\�:u4�(�������}�:k���0}#oL��'��BHC�9}�^�
CDG+�M0 D@�����N������a���ʁ ��p���\���.�W��^dT�R�vjD�5ꉨ�5��]����dwD���]��2��� �rE�(b�6Q15��LdZR,y8g�;�}�}����1�z&ƳP?Uq��I��j$P�0<v�,�Vm�|�a�Jko�\������)q!B��&i��|TC犒�&`W-����[V�	�!�~�lh�\Gr�\)5��{��Ke߀��>�Ul W 9ZM�O��Ƿ��ۆ|Y�(���-Kqr"�dQk���
[OI�2�/�ó�Z)��ŅSx��f��`��X����%L@�b�'h��ڻ)p�߆��R-�ܑ�љF!��M<�a�0'PxX��Qh����ö1�S˙zD�uJ$���?����-ŵmL����,����|�rD�W���Q?�©�z�rJk0�Ci=m�;�<�p�w�O)���r�>��Z-��C�B�3��a�6�k<țĚ�_���ޑ�_=��}e��e���hMa���#/��)�ܷ�J�.��r�H��|8��W^l�3����YҴ���x�|��d���<��0�
�@��a+p5�*]"�g��z��l�RH��]��DVם$���H��IC�����~�ڈ7,,["�{�w��bC�٫6'� Ѩ\�m	u~��R/vN��q�I�(:q:�ײڴ/�,J�H�6+$lW"�X#5�!H�L˄[YG���	ȈI`�� �vW�G�V�7�bD�m4����L{���� �Ŕ)�ݜ�iq�
�+N��ͶZ_T:����ǌ���H&Ť
l����^�|���$� ]��}=Z����^���.����;E+s�]d5����ۢ'�Ya�I�!A�BS���y:���f�'Rwj�Tcq���������!%kL�#O�VK���4��21R�=�T�)G�l�e�,�𕟶�u�ֺ�[���؈�ɟ>�i�ԋjT'o��J�HO�Q���AG.r�M�|Eo�x*.�CwCk)Or���e堁��7H�+{U���yK,�{��t��9?k��,��ˊ���k�6�c�&�h7�1��L)�"� p �m����t�� ��	��ބ���`]�}�,r�x�;���zG�JW��"p�{��޹�@�v��r��Q�4*_� ���O��f�+C�i�$��n����̋���ű�vL��ٸ0����/�Cu�=��+��>�����[��,I'�KͪZ[B���$'n�&f�C��Q��iV�CD>YB�|�9""�I �zශ�>�0��3��<͆J�i����l��_븦:��(��Y��UzZ��Ilo���9���ub�<�"�!|�$y6��n�
��K欸d�#�j�ڴ�fT��f6���i8~vhM!b
+<H���n�S��]U\�m	��!2}��rx���Ⱦ�4���T^sA
)���}����CN�D�[Ac�33H���'�+��W
LF�#�N���o\Q�KC��q��D~o��Y�h��I��[�-Q��O:��UáE��G,��;�y�6��� �I�#��f��R�htव���ީ���^�oѦd�&���m�zy�ҧ&�W���I�垨h�MD�S\bw;�a�?�Em�� Q���&Qv(*_Q)��.���0Gʰ��O(�<�B����i0�Q��)O��"c�wN(_$x>�!��(%�i�|�~���X��`i�!|	��R0��-C�e��+�� (F�C%E��!B��v��2�坒�O�� ُ�	���n!�4d�!�_{�C��Oy�̦"ѵ@��Qt���+�߼D�C}_3�N�����(���\����D7��Mf_˽���� �U,��U6N��7n�H\F}k���y�)]z'F���}�+ʷ���	i�	n�0D�W/���k�4u>���N+��]�l ��9����"o	\�z3_ͪ��	XJ���O�x�/G=u��x%Ԓ�%��ּo�l0*�d�o�Q ��OJ�����X��~���E-����a�+Ϯj�5�:�alEA�р����=h}�cS��0��j���|�2ɨV���!1ߤ�FP�VE���&3���R.ÉDP~dr�U�S>�6o�v�ư5 ٿhe��),}H?��?��1G%����?����F��sa5Z�!F�� y����%r߁%�a<*{�I6{h�n�`(�Q�=�9l>TM,�u��ĝ��2��h{c���w�r�
��`�A�
uq�S<���Y'm ����K�5�Xy�H�
Ⱦ� 6�?`#�1�C�)|CW�ѵ�`�(���k��O�@gi�Ly�z�9�]�¢.��@%)�&8(��Lf�Tv�������AN�>w�p3��������&�6��)�/	%�ވ�pM~
͘��U��u6�7�x��}0�#�)�5]}vy�8Fnd�c{�в�����r���:�3���pġvy���O�U>,��Gj�wM�S?�u3�@�O��҇�6}@jx�lT�x#� ( �Th�LP�����z��
�Ji�UP�@�WC��	�D�����y���]�{U�g�,� "�w&�{��`Y�;�#D��U��z�Z\�|#������p���A�%v3���8� ������&��oY�5�Hq�_�"#^��S�9�����_}��Z6�gJ!��c�_�\^���H"����-�`WU��9�&ڦS��< l���{[s����j,�FI�\܃#]!�Ղ���h�{�;���H~;�+�J�޽�_=�{��NġP�rGsz��1{��E��.����w��-�:���K� �WH��\�S��?M�q��md]Y�O>4h�.?��XS���J� ��\��� � �Q�5,:eK�6[D��"���(�'Ш`ߡ�39S$ՒR��#e�Q�]�T���Z���3@O�ASϝ�8h���֟{f)p��j$��=��:�Uw��i��EV�h���oH+`' |e¼���U�_(c=��r�V�'���6�4T�e~00;�0:�f�C�&l��P��>��I��(��?�/aQ� ��΄f�c��D)^џJ��p�n��"�ނX����͚���;z.d�ç��
�L�7Ӓ���\�Xc�e>Ã�-+�;�S�����#�2�� ��3=�;6|}� B4��;���tw4�7�Z64Ěb���'u�LS��O1F�֡�y��������J9&K����;��f���S��=`G�	�2����1��C�0��������;4R�ɠ���DFK�oV\#0���橽���bu��q��y�� ��c�{��N��%��3w���	�F2�022t�@�Y>����ẫPݚ�B�~T��8�u*���������(���!���K@мG�7|S�%"x5����������KD��TA��Z�0��.ܠ�۬s��{-t��RB����� �N�A�wb���ܑ�6�C6��3�!��t
�|R�b��bj��p�G�����h�6A������#ZZEG�&��9�gU� \�$$�I��O�lWϡ�J���J�,6�v8>G �}�B�a���mL)�P<�	9�`�mJK)�.-CFd�Y�4����ӌsRG����녽Jm��#��Wn�����:J���U�v0�A��ژ��p��|ՇmE/0n���w̛�����'mo�P�q78���~�u�#Gn��L���$�q���ܭq�}��*�*�F��K�2%�NU5�SOu	Q��� 7�r��pa��ő>K �l��CZ�R )^|L>͓},>����j���C2�۞�5���0�Q�8ʶ��I@p��W����bm:4�,����f��=�1�R��\��͖�9��[�J�)�ir���֣�/�jN�Ȓ}("ɨL�8���A���,�~��I��J��	����N�rM;�[8`���C��p�D�	�)iTdt�z�:∰S ��5�&��7�'��kT�ӆ�L�y�'�?i�-��I���uT�̌s�0ϣO�()l,�������Z�e��7*>��I�'���M���d��l��1�4�5H0��1��]:r��!�o�g��:������W��o�'j�@e��"r%�\`J�v�:�ߙ����͑��)ǳ��;)�.}㑴{�]����'y��*�?'4�.�\c�H�1�>�c��N$�|6����^� Lԟa�X��ȫ3�_�3�r�&�A�mbė'����߬@� +9!�BU�\m8%���"��4�QH�/,�2,8O��9P�;V]$V��+����Y��!�C���e׭��ۗAR��t���� G���]��H�}XF�L1t7�G;��;����{�-�_���4��=�J0����ؙ�a��լ�4�)b[��[�O�p13�
�A���(񖶑�x��Îd�#��J(�n�Q7�Zɜ�v�����
�&L����C+�)���*J�yl��c���3*,̮�Mr`���Q�FQ9��U�~�B��O9�=򈊼 w)d{��y幮����#��fd�it�V�Q���5m�L�����H���[�u�uI�xz�b�GaEV��]t����L@�_>eƙ�t	��K!��}�z���R1?��jm�ݼ
��<��.�TN��0G�g�24�L��x6����2�� �އ�S��8��lt1l���l�������skFg���>�F҆�;A%��|zMgmvJv�X���w����S&[e
A�Zc'h)�׶���B�@�&��]�����z\�C��pw@f�Px���DW~q���y���>]�3���9RE崅��0��$�G͐�'�b�l������3�
!�Ϟ��l_`6���q:���#��(A-u��������bV4��"1�n�)[cTr�|aR�0�o�����p!��E%�R��L��:ɉ�Zc���y����}��9�ke�zޒ���S%�Tr
�6��D����Y�qV7�?c�t�R����תiȧ�۰��,�����ӡ�����KG \u�~�Ą,E/灙MT
�߻�R��,|"���$�s���b��֭�<�ƞ��E:�@��M��C�{��g`�T��3i猶&2� :7rUm��?엄������w}�(Yg}SU���zm�U����֯]I=�q�m:��f�'�
F���(�"59D�R��u�h`�B���� ^��M�К�Xu���05Jy�:�emF ke��4�IH�ΟH2�'^~�{_���D��\�d;'K��7�DB���`:S�����+e��g���"mEu�J� ��'q~YqҒH#�3�_����USC���՛z���Gp���DÅ�Qo��>P�7w;lƧ�2���x;��Wҹ�<��.��p�!E�#�,�!y�e�Ϗ	Ou	��J?��D���"�nJ����c��T�e����2�Jϡ�K1�39u��R�3h�����r�am�HY`��r���#�{H+��L�'�j��T陓�Z� rl[����]�}�e*+�D)�����!kWt�?��J�x�]�;��jn�2���S�IA�S+cj���\+���`�vW�ie��,E	"��,�%�5����A�~k�w:�6�h�e����o҃�J}����5��zE��I6��8���jǱ	�==��N�m�
��'��ݷ������:Ȝ������������"���	��4<uC�}�^?t�YW[?W�?=T�Ҷ�����o�wH,����ḻ�oA'�)�΍�kF1_�L�x{�셙H��Xix/F�[��^H����aY#��*��
��<�b:oS�2X1�T/�y�}h����3K��а�q���*J�}=p�eڂ@Y:�_o|�����VuMC�Ԥ�N�T'Óf3�i�\��aZS؟������=�����vK��u|����Ns�� �����5�;;��&2F��Ϯ���ZK��� X[ܜ���pb��=R�+ �]ĩ6�<9��	Q�=�����t*n0���.��	�q���x��ׅ�N�+ȷ\,�]p��ce<��\|�%���AB_oLT}�ᏃN:�C�&;#Ю�ղ�U��i�0T����P3:����N�40�Q`�T�-c���۹�M�٠�F>s�РUaz���"��oai��Gßホ ��Q�P����T�[�)@���5����b��BfD��w�$���o�Դ����)�2���9�3��l��f�yQ��zbE&YĴ"!`J��-���^��L�8")Y��[���9&ҽ���y��0L�OG�������HR2���ݾv�͹�Z�B�K��2_ȴZ�aKH���A�&�zVӱ.5���	s���W�c$$��ܚ��a���g��P�i�)[=�()���r�p)/��J����A^���m+e@4��{������N9�F�i�Xb����pxIO��1�|���Z���'THr�����t�ʸ��O$�Foŕ�m7 �WDH/Vſ��e��KEn�l�H͇���R�aރ6������l�7��H�D��d�C�C�D�$w�f�lk��|��أ��(�������t �<Fy���X��aY(�� ���QFjM$�WZ�Gso9��O�QC�3��β�D(muj���bZ���#Ɍ@�p�;�hp��#�'Y
��ҵG�$�~CWY:p�Hj�v�hH)yl�Dp���զ3z!�����}�SN������B�-��WʖP�k�Zۊ	���qȧ��\�G�b�o a_��'�g=�HGk d}Nf�lXL��K;���Ǣ�Z��eo����-��[�����v�R
�I����/�Qy�Ig=6��4Ek��x@�1]�ͅf�A@k�Sx��յ��I����X��׀���3�k��-�as��o-M^jY9�u+H;=��&�y��k�4ȕ ��E8�D��?�xP���Y�%�8�VOk�)1MF������"Ǆ*pEC����J #�G���`����(��p|����̹<YF�8��:�q���Jm6��)\�J�њnY�zY8�U�aK�s���,x:N�i��a2\��.h31M1��c�<�����Ѧ(80|� $�	a��U4�������͖)L�g]�wo����y)�n�n��+=�_��oCy~rę�3����k�@�d�6�&��+[\��#�)Q�_���d�MQ�2�Q�Bt�!��b���>�|Q��w�2�z��'jz���/��Z���B\ŇD B)�K떲���moâ�0|	��s�5��ƿ	�e*Udj^.��ѝ�Z�8 ��Y��d��F�e��-��0���n.k&�>D��P��ڪBm� �\���*_�����sL#����~��)�����{��l9u)%!�"�i�B��[�
�L�h�6M����L�E�_���
�u'���[���;aT��?D���4F�^6���������838�m�1�+x��|��#�A!�ϡ��t��`����伏�l�Y��-]bQ,�c�o��g:�/�o&2�e8�Q9�gȊ��6]�6���i����0>/�K�eo�+�a�������O��}���2���%�cGO����[�ѿ�h����o⒍�?a�)"y+Φ���l_����\��U�Y�hb��� J�.�'��4��ŪA�σ.oa�Kˣ[���J��v5�sx�W������|3��?;Q?ܝ�\"�jsʕC�%58����9���+ų�[��O�?�ƒv�w2(��(�h������͞z0ԥvU+���0�"`L�'_Ҝ=XU�a6�`��,�H���(�1#4��@���\������aL�
�JC����yVBL��W�	������1�;M	��<��wۤC��/zi�0�.{��ΰ����[?�)�JJh��ɀ)(�/)fNKÄ������M9����툤���Cj����5c�'�3Ҫ-������ס��H�g��ҫ����V%������ژ5�����v�`�V��TEօ%��NN�\��5CV�in�-4F�My��H��{���:����������5'H��&j
h��9B}��
���l9xM2�(�(�ҁ��K+".j�q��Q|����u?0���_�rA�o� �=��B�~�!hd��qa�ۇ�Ե�\0��Ğ�;(Z��zߝ�5�ٸ�)�x��MTR��ɿ������c������ϱ�P�=�f��u�)&���q�xG��� <����4�g]��r�gEfE	Ǥ�6
3�1F	�  ��loZ��;XS�$pH.�#�"xH�v�ǹ_՘#N77��7&��)?盤wl��J.�V�'�hn͂�W!����4j�	\̢�]�6vQ��=���`"�C[��B���;�lo�p/s�����'I���57p��t����