��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%���!�h�^h�Ʋ����8L,n���j-�.��$'4@��*��9�2`cv��o��6����� N
��{mG��Q�!�j�s6u��\E��+��hA���R<���+R��"g�d�����*=�.�+�L�L9�]ʈ�B[�~�R��ҹy�� 0N,Ɠ$=U��_�W5&֦���%�I����-�}ַo"��z��ʮ>jsi�����N�6C|;u���S�@SQ�"ITP!g&�Q�>�B�8q~�G�ǈ����N)uT��џXd?sy#��� G�ȩySr�~�QN�pg��;MK,�u�PL�[(�N�"d�Q���ܡc�·�WQ
��V��r�T��2��p���v�e<ְ`߬���u���$u���q�)_R�7<>z���F}�c��N[q��˖�Ng�s0�))��4�W�x�MO'��)0uE��T`��t�KT۾X����.7 ��Ͱ��E'_^:�����:e�9�j�yX�g���)ш�ӯ���Hy��!��ӻ�e2锚��R������&��\,Qc;��P~���QNc��ty���'�����*�di?�'�@a���%gis_l���jφ�PI�OE�����"�3�$ttum@?���E��w�rf��5^�&!"C��~�>l�H�5���ʶ/���|I�� �l�L�쉯��5$�[�����g*^ôDF���������	7��O6[��Gl2&�=FdқH�.3�&Ȏ^߀�㈂ŵ̵�R�����A���"�W��ܩ��aV�/��%�cl����i�o�R���a�	Y��!l��ѽuS���^�-E���H4)%���#�T�Q��l:��˲���f�oˡ���	L@	;�a�,�����R�z�E�\�E)g_�������`�dJP���R�rg:���A;&�"�X��\������J�B��kF��'([�(^?fo��TΑ֩����	�A8z�<�:~bz��}*7�]Y�=�A���}�C\�C���Y�M�v)6hM�l�D����f9`���|�!��Y�;ｔu��@�����i=���2��|"ם��P{ɸ$[?}�O�T����޼0��M�8؈�1o�q6�(�(��ק�B��UV���\J�lW���n��R�(�����ly��kN�����^�ZPD��I�p%Q�ѝ*{��=w�E?�3H�)�{~p�]>]����2��4b?�mz���:�*�	U��΄Z"+�}�ε��M��!f4����M���LFf�W�1XD��f�~��=�oC��������������k��D��/��*Fg�U3�=�@�NMf����,$t��������P_AʓpH|��|�Ѷ�9 �4Pg\ia/zN�_�F����X%���ۖ���{�^~�N��Z�\\r�j�D�F�kKx$\"uG�G_�B#1���+f��>N�h�쏎"nn�ewm/T��XsЕ�2N�2`��s������#_oQ��1��;��	l���d������X_
�W��~��?�h��.��(4�Jի��n�ߐ���{)D4��eTE�]�r�I�X�L��G��$����urݐ�zO�?���J��L&����ʠ��u�&� 0���b�R�L�r��b�z��ZQb��@vc^�)�� �}O֧q��9|.��"t���g���8ΐ;�D��e��[C��Jx�7��6���я�n򚖵0-���Et� �=oW�haiE�%����pڈA��#�WNC[�K�F�Ow�^P���pm�⼜��i�Fu�L�������b<��3}�u8�+���a���v��2�c�{9>�,eq3y�#u6\���i��eq9u9�C"����V8a5��)�t��j���S� ��2����@M�-B��Ȕ�z�4��.l�0`��曺�L|+u4o�,i/ȭ�Wt�G������7IF�K���1k'��f�zÇ�x׻s�{{s�.���k^S��Dn��Mo�p�X_�RU �C��g�T2�#��X����J$:Λ�qU����u��-GF_5=)�аyM.�Bv������9�֖�of��>~��U�(N���ң�T(��QU��ة�"��	
�j���/  MMU~i�{��8;[/y��T�����( ��&l"��4��c�3�#��(H樓K�/wT��_�g�]8�[��T�����4lՇ�3ؗ��	^lӱ����ٮ�9���T=-��>��A��|ihtj���eO��F�`Q�۶\V�萧��P�쭰t�ynJ��&�>�P��,}.�ʬ�	=x:��̈�k:�k��q9q���@�:kr��1ޣ����
�14�rd�-����\�ԇo	e`��_q���S�	FŘ�*?��l5N�_���BC4�g\�9+H:�L{��vU_G�t�T���bJ`��P����&�!)"��r�+�O�d�;~��={���On��j�Zwa�XB3q�u��Ʈ�
�u���V����ר՗�.��C]!���oL�'�ĥb�[%�?贷%��D;d8W��ɧlj�D�>(r@3�ۄ3���$�@Ů h�7��M�N������F��u��y�}��������ߺ>l1C$��*����V�.���I�B��!����4�b��|����L� ���X�E�fZI��G ���{����1D��F�"��û̚��+
�iY�;����p3`����7�;|j��3e�K���5�a�	׷[2Bm��a�Fc$�p.�"�8x����t-�`�fO�vo�)A�Zر�>6�!���{{>���
��*��k/&=3-+�=($�OW��2��D�zWg�qb��irE��}A�Cv܀��m��M��m
*9l'z/ gZneӃZ9n_-���l��;]���7�B���Q]���-����Iz��h}�@�5���$'5�����X��+�@�A!����2��{
�@@7��2�����D#���*����.N�Ը�s-DBP���٫�6ٔ@�{��W`�Q�;9�f6�Z�1�OW7��9�LĔ�:��#OЋ�/�fMA Z��>����.����+Z�m����uT���y����̪q�h㨲��є٧�ܿ�Y{̣ė;hA��kd`�xֱX���N�`E��C}� W�u���M�U����؀�����_S���d�4�*�ʰO��l�M��RSo���'9�<)��F��i�T"��JP���1v4o�%�����&�e�z6V��F�0���|����|k�RP��G��i�4V��nBl,Z^j�Ag=�$u�sd�+�	���C�؆.}
ph�|��#���fU�Fj�Q����XU'�`@�6.�n����]����-=.ѵ�wȦ�&��祧�6�3����؏8j����g7��{��a+^u� ������Ba��٬�J�pc:s��W������	��$H푹��f���&�R����{�0eY�c�B�>J^ѝ^+���!��д.!% ^Ƌ�6����-�ь$���b��}�T("i��M�B�&�-�������Gr��L�����4�?s[�Jpe5���+@i?-��"�w�>I��>��d�L��̚�җ)�9��*�7t�(��n�PN��S�o7��/�E0l:{��	��9���1?�������lc'�@n��*���f�� � ������)�@����������W����_�އ{N�W��J��3�����>�nf����'ix;��g�6̴�X�0�<��Q	�ut3��\C�ԫ�6�����d$�n��Jɡ�@T<	�_ -o/��#+�Q�=�H;w���b`������GoL�Wz������^��Q_8��e��}�Qܩ�nU�9p�����U�t�����b[�HӴ����x	XT@[7,�3L"���Ju���A�M#>�u8�i�=IgD�-L|����i9-a�%��?�C�E�UI�;���.�oQ�&�F �.�zg4�x��<�IȒ��~>�`c�Ϣ�<gw�l��Wژ�[�k�ÿ�Vnܶk����'�e *���Ԡ4h��Uh�k�W���D���L/Ѓ|�P�;k�D��V}]�Fx�fJ
�4�Z�f�=���E@��_�F&�)�[���E������Rw�H��Mi�L���9�`����D5�׉̮�B�2pK�&"�ڰ���7:����M-2wK-$/��I��+y���|�	iṸ�-��������rlx��1����)%�t@]F���hMF�	r�����k��J�w�u���+9V�`UC�'g���EJ+��n�[�-�Ѻ�۪&�i_e�n�b;�7�юYn�m	[����(~��o��9"`)�.��1�5���F pr�+�l#DG��/�Z]�QӘ��ޕ&X��bĴA���*}et��S��D'�K��/ֆ{WIe��|`(Z;�k�Q�F.��Fq���+0���'��I(�{�rtC�Lz����,ƵҊ��%<��?P���`V�o�E������x�7���?I,|�N=�#�qU�TuI�%���p����o����s ������6P��[�Q�.p�U�Ó�/F,��]�lt	��I&~u�'�3d@�7#/F9�+d5j݊]l�b�����[����r�n�(�����8�Bw�R��������uk[�ѻt�T�@@�{��,��Ϡ��;7����&C������`��HG:z��>�0��̒�'�����h��}�	Z}��������	S~l9���ޏG�L�htF�s�S�������b3�P��)y���=��Br�ͣco���Tz�0#�@C�_��{��DyFq��`ݵe��w�f���5���!�zPbM15��J�N�m)Y8S��qi�â|����$E����U}ʣpMci��-~o|N�9N��w�)D�`�k�v^��Ch���g��ش@ r���;pĉ�ռ2@�fN��[�=�c��/��%V�[�>���w%a��y�h T?n�.`�p�8؍�V� �"g\�6�a����]u��ه#�ݑ�1Ӻ�ZzQ]F������P�KL%O������@����1;���\��:��k�f��V��|�es;o�h%K�����3���TP]��b�� �h��=��1����O���T��8<�ge!A�w��]E�0�����<�=(]���C7�@l�&�����2e~��an���~����[�����*��8�1�O���6Vi# ˝��-Ir���r��q��
G��/��)|���`|%�����=��6��Uɞ��_,[E����*:ֳ�^L��^�O 5o��wel���C�JJW+����F/�$	MX%(�g�*!��+��;s��{Y��ou��6�)�1ee���.���p��&��V���yo�G��iɬ�[�v�m}�FZ����q�M��������F ��Ŏ1�h��I�����Y��%g�<Kµq]�d�����������3��l<>?~"r�^+Y�
;P��_�r�)D��:�����LD�VCY\�y��-.����[LW�&F���F��@��Ѡ&���$�tuۙ���fB�	����<���A�^ծ����7	]!�:ȫ�0���/FI�}E��QeB.��أ�������;�J9�'l��f{�ϳ���
�8V�0��\h��{7&���9C�Z�h2���O����sr8ny����م~
u�!���)��<�Pc��E�n�C��r�[+a��bA,��%�jJ���������e{Žϒ����5#�Uq��kɄ��`�a�!�u���{�(wn@��Je�p#?ಸ�c�|�M|��P���lo��6a&�O�i#9�s��Wfjp�d́肖�X�(ٯgp�֮ɠ̞�~�@����+��ދ'?��Wq�/Q{�;��N��� �(+Om�W0�T�Q��2P�:�)HRH�U��Q���z�qN�o��x�'�w���x6D�S�]�l�Ra27l��s��H�2�<u��Z&���Ixzs�0V�I���:�A�=�@�Y�Reb���f1��EmJb�9��SVLP���$pfF?H������$�Uu��3Q�&ň���w���S�hɅ$����~��v�$1�O�a��d���?�V<3��(��߹�����yA2���9�����8"l�I��}����,�������Nb�O<�;'^�3D��y��r��!�r#t}V��:?�l�hR�fʱ�JxH�j؎��d��c-��j>��~v�{!łXU>���1�b�Uβ����E�c��jI2i��z���襝1�c�P^��� �5�y�`�$p�!� ܈n�Q����[Z]A#����c��zC��n�S~����
��շ�J�<4x~�P�����#F���Y���l�h�q`���v��(W�ѱ3f����G}�%QQ�^j>�;��1-��S�ןKN�q�B���sB�>˙���[M<�?��E-����¸]��6�z�ȣ,���� ���������2N݄��a��lx�>N׋����1�Ԓ��lw脥��4.Aʝ�l����N���	ؗ�'���IS-���c�Կ�;f��tQ�4�-�ڤ|�Rq�^��֋��b��`��ً�i`Q�cL�?�Y�)z�0C�9�rp�a��<����A����7�]���Vς�nO,��f_V���竴���f���f�e���0�]V��97u���fWK�o�o��R�����򮴕8%�wD�q�þ�j�8I�m�tUmd~��kBR�F&6*������3b �����3�6�-aa�kw{����x��ƚc-�.Dv�->�s�w�&eLy��)�G�$��X�_�_/����}]J%�Udr1R��T�=�o�D��{hl%��q]R��Wy<�s1�ϳf�
�.e^�է���	Ҝ�(+&�r`�'܁�^T�C7h`ܴ�寲�Y���(���i��gώ�H�������H�v3QA��/_���