��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��׶8۞�@�\ږwiܕÜ��=r(ro�fC�pr�L�O�q����6�|��3�Y�	��9t�1�HKjQif,br��<J��0����p�l�i��Z���T�Oׇd����e�/���x�\����l��1���F�.�a�f0!�:�m�y2���u�%R�k�a*7D�dJ=��4���W�À0���2$�*���������v��1]a��oB~L��?H�߷NO��uC%�h���!2�У������$�Q�4�F[�2�}S{����$B_�~g��l��LlQ�tA�|��箿G"�M�xk�3�'@��V�ҵi� |V�(��1����7w�x������0n���7�uy�-�>���YG����￤-�Z��F|�.�F�F���6i9���w2�{���L��RCj�!,J�n���v��*BOV�*��B2��Wf,�"i5ᶶ��i�����;��Mūɝ�qfڀ�-��-�N����=Hƅ�ǭ�
U������$���Ǆ��L����H�8Kᾚ�V��E��bP�y�"�gC�塬03����=/���ZoX'稿A�����=z�*ì��a/�9�iJK`�9��՟~��F�נ��
���JXM?�<���Sa=ǃ�# �Y	L���GI?��D%v�^}�����(��$+��Gg2�2�1 ڮ�U�Wy�-��-c՝�BQʎcE�E���+����h�W8j��G$�U�M)�r�Bc�������T��]zBS�;��-���sW)��ی�!ַ��=4c1��)Nf�0�H���<$ty"V�a�}��{���?�±�+!�6������">����)l�T3LeT�l����5��߭(٧�4 ^�ţ�(��ҿq��]>�TԿ��Z;�h6o8U4Ō��niKu�i�.����#�C]��l��k"9�j~n��^��W���O��x"�hki�߬wx�.[>:b;u�g���ኊ!�{�Jt"����o�V䃼)xӀ�gsQ�.��?s3�`����M�1N>m��
,��g�d�s��f/�ЋŠ77Ξx��� ���6�@�8�-�趢-R�~Ӡ�o�w�P�6CC�a�7fߪ��'�=$鲨��Y���}:^,��<��v�]��֕/� ������:�˒���Y�m�&׹.�Yc(��ד�p(f�7m;�/�7ch]�.�K���7��}$�pr�"X=sCQ�rB�y�WL�_-H���Ii8�AL iе���ݿi����m���\M+��Q�O��3_�.�#��w�As�O_�V)͍et�d��G�Sap��܏rv»�7KѦ�if�VGp����h�$^�|̘�f�� ��.��' t� ���I�"��R3���Ò��xB�^��VZ�d���>�A�Y1���1��qX�&ӶH��"U�el�d�c�����X)'l{�[>B�M,��ö������M���5�����f���
U�f�)�1#��d�:�3($w(������Q�Ђx<�F��������#�U�'qS��� CK�3p�w�4]���l���cBi�</8�
�(!��tV�W*e���^�L]`9�[�(7��R{�u�b�-�8�y\���kPCR��� =X�H�ڂHt�$��f=!6X�D��Ζ�S�+���B,rr.ջ�D�Z�C�+�B��M�T��q������oR��=��#�E[�P��h����w��j˴6��1������i,(��62����'�~��[����{#5��w��ͦg�3���@�K�Մ"QZ�7+��i�Җ�H�"ϴ�gq�~�_(1�ח�]�r�7��sl��	ժ��1!��P�ƺԩM�{ͅc�MDq����ڳ�xv4Mh���
��xB{���	�d����&a���1^�dX#It�w�!���̫���z�����jw�畹��{@�������ϵ|'o��cJ�8��NL{�r̬NZ!�a�ϫ3&����jI �Gi$�'�� DGl��5�}~���4M7��3�l���_-pG����gL�G�"��R��|�3��\�$��Ab���}��9�mb����{F�t-~���C'��A;2_�R,"�@ �^Z|ZQ>5%�m�j	!F�IR�`�Z�E9��r6��H������\���q��M�m��y!��<��a������E�ކ��7���&�6���d˙cv�v�J������k;}D@�*�L���lH��M�l��Z3Óz7բP��㤹3�-t\�	��f}рt�q��ڨ�d�j�J�.\���z'���.�1�O2��9�ѻ�i}�1�vo�
q�����5���o�eh�w�G"O&!zl�ϙgC;��wz����T��*�8uM��-�8#��(ͧ�nBzH�)ܟ�p�	��)��EM����e��	ї�d�@�)|r��޾ϒ���6����Ƹ��a����۫F�.t���:a�mY���<&��]���L�$B�S�Mf�?qS�z6ׅ����G��_��-�e &�q�,I���`0�Xۺ���y�QH�^'9ʞ��ց��X_|�i�W ъ�\�<�+t�
%BP���!�˃h�j@/�pi4�"�Me4������QA�niP��8��ʮq�Dh�+�;{hƜ_�����Y.&�ku��:w�'N\�`(�w{ɲŊ�G����s߫�u��=��Y�`�����t�,�m܀U���Z�� �i�T:W��s��T��O9&�����z"���˪I�˔��ՁIw�����۴9< 80Z�0�x�zc͢h��y�F��1�k ���Q_؉�#K���L2��J���#3��)2�m���B���+ə����M +^'�1��I���d�`�1f�Tà&a�)�T^:\P��A�cn?Uo�]�s����nmb
f�o����,��Fq��s��~��l����x)� �3}X�}�^M&5{���K;0��C��/b(�GnZ��#�ٴ6�WJ��6b��n֡��|FP���:UP��e�p�Y�)#!Q"�7��T��/��X��ɉ��$�P�Ѿ���߱$�aM�2n��Y)���.�a@Y�������U�s�c:i����T��b�ͬ��X�3��FF4���ƠLR;q��]��*K�9��2���7��E�����mi��/S�_�ŀ+Ύ��A���v�H��tFV#?k�g��4L�3 �2�N{hXXD�K��B�-u��e�5�x%���cޥ�.���n�9׏�w�&;� ��ӫ��H^�w�������AN�����x	��F��?�Ƈ��;tDn]�jBO�v-��OxmX�6CB&�o�Y�N�q��c޽[��Z�M���� ~}�ߌ=��'�'��+C 7h6l0��f'IΔfi&�pWrv����Ǐ���/�&�'�ɇd�2���I�q�>E��|���Cd����p��>,�plG��`�ppT�6�|>������R��B�����	M��oQ��j������P��J?+t֘���A�G
Վ-�o���I��yh��	]I���Z2&�}8�Ɍn�|�L��Р�6Ո�������߹�(��N"��6��ӎ?�E�Q�0v<�V��Ҕ����h{�x0Q��"��v��ei�tl�3Ҧ�(��!"?
wp�NA���C���!W�|,�Ԃ�ٖT�x��y2�n�>{Lb�X�3�:��>�V����*4�A���:�i���r��ҳ��yfį+2��T��+Z۩uIZ>�ݳ?a���ˊ�*���3�E��?��ʯ���k�cC\&�
��6��z|v<Wl�s�
|�����^�'��Dm�@͆�����0�ɣ�͕`�21�_�YXЖ��i���{�&��g����Y>su�=�59Ҹx�m_h�£z��nm�3��2�X�/V�Ύ*�|�mK�D"�կ�B�E)�g����&�m1:��T��h D���E�6$��1���ʠ�)ϼ5��W����8��;Iտ�A���?��]�pB����_|Y1��r��JS��E�9�����c�!��)x��o��!f���[�_�w�3h�We�u��h�s�G�k��x6�8~�?��u�ݥϰ���h��}��{���^��;���w�8IK��
�[L���3��^��>�2�oQ+*F.���4:�oܵ���[<���Uڵ�gF�A��$�^4�����$������<�Y�1(6�ۀ�1N�P��4������� D�J��Z�0nȣ�2a�qe� .�µ�m��i�9�ܺ�/��W]���T������ژ#�6]6P����30?s�Iv؂8�·�(��Hc:�/�,�edz�Z�~���Ґ�	��N��-zL*���Ry@1�(��`�1�d���!�uae曂7Ǎ�|�D�u��F�0�H4:����C��@�Is�<��B?;A>.���[D���� 	a���`B�)�K�y٩�
��+�6?:ۮ���P%_*O�J�0�����1�+���g��w��o��(P̨�6��hDb��kb�)褊ʗ���?�L)o��Ny�ƄA�N�t�bW�}^zGkj��SHL�H��$�r�a ��?L�G��H���9V�n�ZC g�k
|\�v	�ϝ�"غ���n��g�M)B3�Ʊ���sc�F�|[��6��O�	[��[徰�����	�y��u҇2�ۚ��|+^֓���:�c 
O��j�{<��cm��:�҆ $�w%�L"��a�/��,�'�K����MÜ��s6�<D��7')�"�.1���S�۹�/�9H\¨܆��u��(��J/Qƹhȕ�R5$⩞t֮sr(ԖV�~2Y*y����ˇ�?
��+"쨹�J���鶮U$�l��4���nԆ/߆��L�=�r��:#Z{V�Қ:����eȫdnr�:�1`�D�f	SZe�nsUv:I���24�2˽�uTbR!��E@�n���~�L	Ŧh[�z�en`e�G]�����~ݓ�@�{� ���/��b�|�y�_�8
)j�`�T��a�rG��,�O$�Ѝ
�o��TNQD �䘐�^�о5fl��攲E�1��,ݤ  5 �U�Pj�o�p�Ry����#5�X�؀�,W����d
������^HZ�A\C�8;�-G�0�_?>�1�޳|�Ǝ�^-x�į)
nr��P,����a��.��@�WE�D�X���VZ�،�.�[]:�`���.��{c	����,Kw�(�� ���3`�1. �c6��+�*�3.�{h�&�C���<��(o�y#���Ȁay�$N[}��@S(�$�*�n�=i�4��T��%�U 4���U��l(�5��;�}�K� �����\<v��B�"Mhf��@�hI(�|�L�H[2��ֹ��@��1˥'�ͩ0i�r�'jVr���v)�i�=���K�Pm��ϓ�.D�{!܏qņ�~1]�e�"��@n`u6k��K��|�ql���c��¿ªR���͸�T�m������
~��f���������KY��%u�΋����ܢ=�wZI�As9�(�0�#O����웤����)fqX���H�ū���!�'I���t������Z�Y���A��IA��2X�8�_��ER�/s�B�����$�