��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQH�x�U�'�'D�~�U�:�Jvx6�v�h%i8\����h�D�I���L����J��z��x�`[D�@����n$��e�e�_R"�w��jp�!��n��J���o`����q�`����tɜ��*�c��s�S�ӯ7R�$�*.�|������Vy�>Γr�t���d�9)Ȁ��l�1���f�w���
'΋�Ճ�5�Mt:��Aka�Q���f�_��"Ȳ��Y�q�0;�c~�QVdoI;���5P8����0�c��k����U+T���Ј
��@8d�"���Oˏ)��zD���oY�p�r)��&䠉�~��P���8O��2x����ئ'e��H��/�+����h=Ɵ���"
R��iw��w?��ܫxUH��j��m:�3'?�O��S���5���,=^�Z}8`ؙ\1����F���"Yg?&@�16��ʊJ�\d)�p�	�d [=)�t����x纱���<�u���߬c�e�G�޷��U�\Uo�Pk�� Uϯ�PކCF��'I�U��?[����E����2s����h��/�x�#�&X/Έ:�à�z�<pF�1�]������ѪHM�w�Vb�K�Y" ���i��zx0F0!]�"��1��}&���yp��R;��5�Qt)�@�V*����4A��h����Z�^$��G��Q����>7�g�@$΍�^�;ri]Br����Q���pY����y=��R�\z�Mmb�qp.�X�X����#3��ݥ�M�V�Y�yk>H�΁�{�c���y�o��u.s	��<�7~0��@	��+��&ߺ�P�.\"���pjM%U��ƛ`>7�3����Q�׃
��B"���b��`�gߵ"ʘ�H�b<yA�
����A�����9�4��{'L>Xh����Q�D�ݕ|F]U�8U=��~L����?�n�Wd4;-��Y�����3ӔMSg������0�X :���
V�Lg��>������ګ�a4F�M�RK�9Q ~9� �l�HY��W��ϯq����6���O� #�ދ;+@u��P���f�`[��1.��/oI:1u���!��l���P��W���ۘ�n��󨁽X~����Q����c�^�����Fү	��a��O�Ѧ�:�>l����K�K]�`�'y�kI-r�8���F�C�F��E�4�ꛆ*���E���L��)4A�d=,ix`j��h���ر���e^0s>�d�t�/� �|Kp����U4!k���&�3�m���,l/��8�t$㻃�/�&�үږ��,fn���(9 ��e�]��iw��Jk�}��c5�Νi��M�X�!��R��Eh�����?1*����`�+z*����:��(l7s0u��l	����ʖ����8�K�
��P$l-c~�O��k���������+
���9?uW B�������O�0Z� $H�0G),���������e�V���舄����Jf���t��ik��s��2���,��rY}���%CRt8��p� 4��,�q��1�R�]��	�`�R���g�B��~Uz�����w����;	4�ĺc�%]&v�%���~��]�* .�Y��8{��/�t��pju����P���ņZx�>_�|�a��0L�R	����éo�A]n&�c62H%jD.��0k�4�G��ƬB �Ղ����pc���(v�D�aN~t�t�"e�J&ą*��ൾ����5���:AJ�"���W@�u_�1�gV�x"�gV?�~�$�4��Y4k(���Z�Qd�]�v�ٷ^�]���+J��tF2��n� ��_L>F6�ա�Y�ð5k5��;2�2�4�q���\�)�8�
B��&Q6��ΰ3��簞U��u?��!۹h;���ڭi�
�[��
'm�@���w�| �4KFa��5�Mہu�-���ݴ��H �j��c��Q���/�Y�b�cM(�,�L�:X�rI�O�`��ݝM ڰs�F�;�� V���ֶ9W�5F6�Z���>Zl�I�;��	˦
�#���wxQj��^�^�\�/(�s���X��@�Zv�K��Ҙ��{6��[����!%4/,_��OjTk��J�TX�s<�RR�N��j-9e�Z�#h�G��P�<�VL4~��]L���O+k�����.��M��5Σ�uЮ�{B"U��a��z����iX�ajv�����"�(��5���i�;T_�-�#�|�2c��1uCw{��$���B��%��B��,?����I���6���h���8H��HC��(�������4r�86
���m"K�#����t�[P$��P836�G^���W�Q�~�Ah8��>�i> ٽ�����/��T�Z�}ܧk�)��S(X0���kZ[��'Yc�?�C{���������ƀ�[؋��g�%��f��>�l��;5����� P�?��~�?zC���K��J���cE$��.�-)�BT`en�Ŷ�t;�ݚf��I������6��@���"�ᱸP~�u�ػ��n�m\��h`�U�	a����x�Z�9?$SE˽��Ȥ1����5ISQz�B�*p0�` H^~���@���w���C���!�|OE�6.�X��*O�鉣�J�C�SU��"����Фv�����
;ZR�������z}�Bo�3��K�/��ӻ}�Ea�R�Cr��%���ɁV��YN�b�.��?yE]%Q�S'�!g�xGY��̹P~']8Oѝ�Xn%W�o����;2�4
��T�S kC[.�����,<�?)6�8v�s*R�b��6|�q�#_b���S��ڣ�[y?gp��x�+5"�
��0��|I�h^��٣n�a[3d��F{'Rj��v#MnF�,r��*~�EKp�3�B�_.$j:�ԣ�WL�*�z(�e�UD�|��*��� ��Wo e�]���X�P��.)��e���M�ԧT07A�G"ZaCG\/�;�B!P�u����h7R�Z��,>Zb�O����wbH�u�2<�)++�Zͦ��3�X��!�I�� |��މb�0�ϧ�K��T�X�DP��W!�2M�8�T���r�j���n�Ph̡l�_K� ָʖ.`��3,���:��Z���p�w������5p!�+J���X�+�*���mC���sX���G��7km�u�0~��h��P�^��m߮
IPT��l��9��ZQ����r{8zf�.�ғ�Q�QP��o��ړ�"����˓��5��q�l��c�0q�o��-���S�ե|��SZ��;�������y��B'L9x�|:gpt.���vO�,j�˰�e��ߧ|(J��2�Oy�m��:�P�.�)��Yy���Q�pR�����(fC^�Hh6ҡ��~Z#�I��w>����\)H����+Z�A]k��rl��Sي6�z�py'U�����{��e/Z麗S|Z�ZS1\�홈.e�{1��}�-H�M7ӤFʱ9D���Tq��t�.v��co�~��U�f_�Ħ������t�#�p��9���e�����L�u�'��O���'�T u){B-6��ˌ���ל'P�I��i�JY^qJd�~������#-0ݣ	����O ���E ��ޓ��E"剫s�.�#��k��Mw�������D�	� ��s�m!a��PN�}���_�L�F/��~�����iN�r@Q*��_��6)�@��i�����L��]�HЉ�*Pr�*��QR���E���ݽ?�1���s��R볼�S��ٝT[|n_�o6q��yx�m��:pV��p	�߱#<0~��3Ԕ �;�,�ǔӫ�}8���yU3�$���]�xdT~TZ[�3�9��ʂZ$�׍��m��"^��+�ۚ�m���V�>��0���ru��Y�K?��Oގ�
�聖<�Xc�����7�� ���D�`fH&�'C�㰬�*��|f��o�DT"e|�S����⮛)�a�c�KZ�!^`�(O�<C����[l%�^f�'ຐ���3��m��<d��^�=hIWG�|����!�ޒ����J�[���.[��8����ǎ\Ee�b<W���f�@�s۲m�^��԰�n	uѰ�K�e�(�mW�*�W`�b1��꠻Q�ݘZB��cc���M��Z+��Út�����hM�� �n��V�u�C�z��W�WFD���%�dO�v�B���'����?mS�d�:�`�E�frw�2�z���q' ������YKӬL��Z~��͋�Y����i�˰�W���p��Md?]'��a��ޅ�3��]�;�Iۊ��B@0���C�:�O���H�	yE�j hFM�)-�#�G�^�؉�u��72�{��O���Q��L:��JWd�U�R�&�4�"��#�vI���{Ul�<F;e���Lc|�;���)�P��w���X���i��T>�Թb�7zb2�'Ԫ��� X2	P-�}d����'��4�V�)��]x��	���o�p��c^w0�.�"(�X�F�����C(�b��LtZ�ۆ�،�࿗��������F�$��-�R�\u�9����zk��4?�44�(hu�g�T�e��ҬǈS��?/�O�N-9�-�Ap�M���Z�e�	=q��|�v�3�UQ���v-�8n�[g�8�@U<�&�����_����)����+x�v>����U�ZK%[��/�F
lP�!��(����b��`]�7t��� @Zb�Cd��68���_!��h��� wM���3��/=�O���)&�8
�Q�pz�U�g�z�3/@KO�$x��l�/�^�1���N �P�e�y��/�Ħ� _+�M�A֡y�y�j�Y�/A�*H�gx��Rd��F��A�N6�@e���;W���
"���22�sC��6�IWVc!^��d=?:�e��h��������.�*���Z#�s�ډ�=��#��*�ο��; P���ro���}� UE�:�q5\�3�ތh��=B��'�&_�j��Wm��n:�B�$㜍 �<%%�c"�|���&�P�n$=|{yH0��"������'5,x��D�,$�l����K�\�B�\�4wV:wҖ\��L����ӎu5�P�`U\$tط�ߤ�7�uà%�hh�� �9q�J[{���6��y�R���J�ZmS�������8�$��B�9���r���Z%�;����_���5�b��A��Du"�u�bo:\9p�k_�d�C���9�q��/�� A�9�aH	�{�A���!Οt,ˮ_�j9f*e�?�k�9�������ӑ��
,rX@XL�@���뻈e�ǌ[z���� DI��s��>XF|&nʧ���ܘuPI-�=�e0���8�+W��tE�Ʋ���D�pK(0�?_�|��������L��:������|��l�`���-�R1L�}(�\\�L��%}m�l��yeh�g���Tg��O��Wx��i�q�D��^�mC�3������FFX�T@ @h\�����0�������iE�43�6�@ܗ�����X�YN����we,��7�9�1:;�g�,
?~׮�_>�����8k��(u�s\{���5M5�A�{�c�[>I�Y-zuԆ6괁��D�Z�eF�������E���v���l��C�+��Q�N���4�YG�u�2�̚��&���r��79�5�+�\�.�PIZl�' "ԩNm���� :nNPV���V�h��Q���>�#�f|�c�X*��]@���N��;8�u�h� ��Z-*BC�8?PY�z�m�p��u�� �F1q%���j�U�V�{���״��a� |�2���6��lJ�*;�O��? �2;[�y�z�t�)�`�
���K��t�KH�S��������2%���D�:*����(p��9�1R�eֵ;z�"u����-vz�œ^�{�Gv����4�lg�z�K�9��a�sv�z�f��K}ϲ3�$�}Rc#
������ m-[�%�Q�$_�+�;��"�I�޷�Ssg�y��*�+��׍�PX��i)8�x�c�>	�
}P�ʝ���Jm=r��i�L쁺j���x��h �����x?�5D3�B�>�W���ˑ���͒6�p�7��M�a�ei�߼qu5w�1%�=R���3��Bw/�������r�ft���x^$w�k�dQ�5㼉�JIF�-�� �c3&8s3��9�#��!d�`{	{î[����W���r�g@tgh��ԓ[�f0{�u�{2&<8��t���h�e���x���'��8�!O��
ƕ�%�h�@�$u�X�����(\FI" o.��z�ŧ1�ƾYn�ڐS��?�TXb{��ы�7ɢt�wЂ�fQ�<������?�.��E��yuP�{1���EY_x��Me;��:��@L��j��/0Ni	X�bBW�`{_�.��g�=9טv/�2���d�5�6,*C�|��0��vX�KC�r�����V�$]���#�lY�` �E�`�"�����k�$mN�MQ��ݶy,��=ߥeay�%�$}-���� &��Bc��M�����zT��s$"�m�ov�ksa�H_z%�:�_�b��ZW�w��}MZ*ѨNmב����L�J�+�I;�	�)���EB#,.reP�5r�:r@yB���T<��Xy��֩���7��I���5�V7�V ���~�nS>�:*�b9l�ؐ��og|_R�R�&sq�vc���(��X�"���
�*�:Ucې�L�J��*J���?C��Ϸc��������8V����e��Xw����@r�#O�h�pju!���������p��꺘��S�'���*���}�(ò��Wx4q6�п��S�'�T>X�x線|Y��s�>ڒx�DG��g��#� �n�t�ɢ���FQ:����&��k��� Ў�,� 9�e^ّl�K��Gd�&��P�N���q����
S��Q"�{�ƍ��諦���~�H�n�������OaA	C�E&g,0
���d#�@�0��'de<�8b2�s��0�I�N�\�2]��œ�FUd�6����-�6x�����g��90��B�-�]1edmZ��^54*u)��yn���Od�0ln�)����m�ѧP,5��8X�N9���t���W���Rb�8&��� ڃ�Rr#mb��l:�N:WIe�sj�,��SP�7{Y`�Ն63\�-/�J�P1���[
v�ԑ��j���"��Tp����D����VKv6�؎7�T�����$�ЁFւ�a��i���|[�m1��R(�:6&����pkd�̭SR=�Z�	|gt�KzY#G�5�f���H�M�{zN�h��f���r/�s�@I�K�*�C����<{��C�"g恀���Q��Z��5�K��
�qx�^:�7�Ħ�]�l&U�����Nde5��L�e�|VZ�c�#��&��~l��~c���ևX��<�� M�9C4{�8㔞�j�5��Bѫ ���7��7�"��dcg����+7��"�^�p�㱕�VH�?��Λ���4�D���툦&�M!	>�i1C���F>MO���+-ܛ`�j�!���`e.�V��C�@:�%RJ���F�|��%�=nr�N<�Q,�Zh�z�O���/� �O`2��g�c��� NǨFH��M�7�ИT���c��R�����Ղ�(�S�������.\ۦaq���^�sՀP�l��48!�h[��>a&v���J5�$��w0�q��*���j�T{��t_[���XI`���+ì}_F��Ӈn�Q�F�8[4�s0:��=�7��=��L��G�Q�5?Z5~';�gV�����2��E��㯋ʅ�����x ^aa�#�e����R� ��X߷�����r���c�A�[�-��O����Naq��a�ռ��S߶��ch���Ajs��a�j�d��F��s�S)"Ί7�J�|������|aX�Ѳ6�FhI2�^U�M�ʘ�Z&�L�my_���	�L��vD5�E�����DF�'(n�SP��e��0�b��v܈$[�[�F��'��<7�kr&� ���s9W�d��z+4��L��o��/�x-� �g�J�P@,2�zE�
y A��P�gM"Z�Q���H{�s�"Iv{ƚ���h_�������}(�0e�?&�K�k:���<h@pF؇K���y��[C��U͞�*[�a�Vpu#g� 	�)�s{���ٷ-�u8�82�-ɦ��t�͌��
�s =䒂������T�PA�픑����l��w�d��p�eS�
b�ƺ����ڤLCe��4Il}X:��c��(r�K����Z�~�&J�hކ۝�ft�s�f��9�J[��e,t�&�0#%&�\���l�'�5����P��-�8�Zu�=�2G F,�~�ȇaɯ��eU��n)����c?�\dQ�)z����E�,L'���t1b�����,��ۘ}+y(��ra���+nI�����,�r����$����� rcP�mwZдI/G[�ѯ��(���z�D��5�<�Ϛ�{�^%3/�R �<�<s�W�J���?(iL�����&��i���q	�m+6d|󱃸��]���*5�)\K4���o�;K�ۗ/�x�ɆTx}�P۰�8�ك��'d�Z�*�M�|�y���;
�[�^�K&�vϮ�?dL�b����g���R�Y��?��mb�����Y�M� �1Ԣ�6�k[�Q&�gy���H)(� �ᱲC���4�LU��VP-�l�Ϧ��xA	�k�������c��a�tXH.Ӣ��&G���rZ��a�`�vM_:'�,BH�<@�f�K=sc׺��R��:��]�ןɡk��D�Z��0�%�VŨ<m�Ō�Jh\_��d�!�糲�+�˄2���k�+�C4@m)�:��Pʮ�w̉��3aI��ݚ�i�ݙ�'Kg��-�O%;��|je�o ����hKNo��	��y�C�������^�^��G���+�ŕ�;�lz�aH8�����8s�pR�M&@m"����;�Z2RP��kM�.6�ax��)�p����<zFl�\��~��"�k�c��a��m�[Di2tA�P��b���W�a���."2�m��Rq^u�92#��x�M���`��E�~t�_�� ��X�w]]����f�]�3>B������Ed�>Yy�d� F%�mX�T�����6������:$FɁ
�;�
C&�����$��kG�A�E%�.�D��vߕ�\ܺ�_�B4�Wiė���0�c�0{��>���G�K��ш��CD��6�'tp]G��&��<��H(U�¾�L�7|������y�~�+��yIo�U�>^�Q�w�^Z�O,�����`�^�0ĺ���PA�[�o�!�孜R�T����U:�ݿ�`W�~C��e	΁���]sΝ���P�`��W�H.^���E%b ��o_m�Wn��^�%�Z��y!��I�l�%���SØ�����#���r�ho��]Kt���pd�g8�<��x�DH��\yΞ��+M���}��6�p�.:���֓J��o�%��'鏅����6�6�?��>v��f�L�%�D��r=��oAPBt
9��+h����mXd�t��-��_WT�̈́�Aq�(s ��%����c�6�n���`#�^[S��L���.��wh�!��`7��/)b�ߨE���p��@�P_�Z�����?��<�|�)�읜[y�{T䢷�C�Cs�7�N+\�>4O�4��U��7�ዥ
+��Ǫ�vۄͭ �Ex�7�.R+�hU����Lg�m+PQ(c��l9r��&� %9�=G�_�ρ�L�	�>� ��l�:2s}�c�$�������Xs�Ccӗc+k=�"��Wt�����ځ�mb�=ԝS�z�ޛà��Q��$�p�M)���BG�itp��_Ŋ��<���p�0u��d$�^�Ц��l G'8'��>�h=̥d�F7�v�f�p��m���G�������[�=�ƔܟXu�pn�ɵ:փ���b��D�{��/�t6�=^��yAŶ��'=�oEg}���w�ew~�M��î��\��:���2��
G �[�$	���;C0�)���A���
�q8K�B�B�TW�#���M�S�Q(�b�
�ԅp�nN��+ ��/]$1䆤Z���� 6������������/�T/����>�M)gPc��Y�l����QT��H��ߧR�,jysT>�7��M����~�&8`�U��V*��.߸�E�/��V����"�kxo�����1%uT'yÅ��O���Qh�~q������@�/�YSӿh �N҈Q�w-�:d*�f쯼)Js�a��N
�`D�h�:�r��\ &&�$�Nے�d���ú���6&߽;�W\��b�O�����Xr��F�f$W���4{�|	�r���H����	�Ҹm�B"��T�,��v]�":����c>A�I��?{=Ci�PHA�,� �����֘�?T�C�Zl&A��lo��g#%o�qO\e��\T�9���[��+@��u)��h1�/��7�*��&cߪ|�"� ���kض��m�#��i}Ӡka�!>z��������.�a�i٢Z@�]�@�*K�՗��mV���,��q,@4l3�oy�⼟�7S��y\UzHg�e������\"�=��0�{�$b$'���$U۸6��,�;۱a��-trD���&�z�}�g�wN��[�m��A�L,qx.�%?���26�H���T�3��h�>��'�v�O�AeC	um9f�?Q9e��7�l����C��Mb�W�}�Ns��F�
�Z7Y��2��"u	��c��4�8����8�;��<���:�v/wֆ���Q��� >����#`���iu=�r=�q�S,�)b=\��a5���3�z7R�U"C�&O��P�6B��[4P�nz�ݢk��K��1&������^�{�A�6�kI�͛Z4:�r��/�s��`�r�h\`��.�F�
� ��:,�=�dC�:�
q'�ȕE��3�<ҹ���?>�z��(�_9�䁷c���FI@2�&��O����S�� ݧ�$ծ�F�[�)�y!��`Rk ��%��h�L�[����K�E݊ha����,S���R��)?��J+e���n�`�SY4:[�:�Iu#��'�܄�c��j��R�n�"����7'%i69��}��mb��z�"
�LH�1�7�I�R�����	xB� �x��,z:�cqMְ0�~����;夕�!�}��4V3]��t���J�N{&q�X(���OUo��دEtu�.�2I��w�HeU��.��L=����|q���:�~d&�>S,�ſ��oЯ�tCo�E"�k��<����W5q;v�D<���t*)�׳��jˎ��)O�|��[]������k0��_ee���Ē ��s� �X4����Ye�!6	�g�$A�=-X-�%�{� L?�����-�uZ9Qp�0G�4A�ix�ǈ�N��_D�������E	<Т������7T�<��~ilԑ�{@[ݤ��h�Qq��׈�q�'����'9]wr�bm����5����o���P�TuTY�E��$%� 0Ͼ`����4�I1����<�)L8\"hio��1eh��]}���M<�6.w����ò�� R��_l�[�vv�ZxN&=#�����ҁ����c�g2�;�o�w���x�CPW5ސT��\Q��g�Y���чA�=O�J�%xJw��=����s�B��6bzz#!9oH���"�:@B҄�d�ݔxqQ��ƪ^���"a��D�����M�-:n�r}��du\{�.9�E���AE���S����/_��4q��"���$T)ԲQ+V��s��b�T�M>�Bۏ��s�{��GmAd�_��6fي��q' q��5y��N��z�`�2토A��+Y�@��[o*�.!���!&�W�j�<2Fmו
I^����/�S�2�tҜ�{(���ߥT'`�-�%C�����ׁT��A�l�`2v�;��#L�Q�D5�������P4#���o���ۡ���(}ǩ���$� :��7#5�F�C$���q0��G�wIiR���k@<�7K6UK�4�^-�r��df�|f���:��R����j@*Ɉ��x�D�0@B3*�v�4�. '%������2q6B>RXd�v�_�� ��~��e�dx�PJ�oЦ��ȳ�1���.�(���QyDL��4����c|i �X��E@N��JN��,I���(�>1��W��.��b��i"�ʸ*�?s��6�ndt{^`N ������`����6Kzm�����y[�03��Zg�2)��q�Ė��n@��;�{�$Q������"ͤ@�D%��C�K�ܠ�h�@��M.2��o� ��Y�M�i�1�� ��WJ��&Wiށ�^D�e��Y]�tCs���-P�n i䰐|�0�?\�����������C٤1Nl�q��ǻݔjx����]p��w�	r{��#yct�l�6�M"�̚�)�]��
��P�>���8Rh(��c�����x����шC�s�^���?6��IH([�ϒPՄ�̉Ӄz��:]�Z��B��#�s�G��@"��S�91F0x����<_��贑tCO�� F��&7	��Tߚ[��1HI>6���\}�vC �/V�j!9����:�Viz�Zv�b�,u�P�|�L�����rК˵�+�=J�[e�V����Ɇ?��5�0�C"�]�)E{�.��I� :cTKdg�&�4��Q��z���1��0�7����MY��Me�'v>�ol�uSN鋢�Y �h���X4-�*3�euN����<#/3}�Q�r�XZ|�Ɔ�K���ޭ*����'���
s������)��k��U�]��C�k��R+ah�ř��r�Z��+�"`������|�'���OQ�34���.�_rB����!pf��W:��H ����r۾Y�*[�!&wʏ��52��0q��ƁBT*8#M��5U�k!�B�?��M����ie���.R�{\���s�����_�r˴7/eT��%��)�t�e5g�����8L��xZ��Ɛsk=e`8-��ģ�e�z���I���.X�U��`í�+y*6+�lc'���-/��z��" 4Ϡ������q��*�{V0  �h9ȶ��"�<�촇Bk��AG:K>��� N�v����0j�&.xg
�x<M�J-�WΰlX�	2�t{��zJgE1:hY>p�?����92�놀���lg\/ u��}6�u_ȓ�Yi�m+�ٱ�	���2�=�±��g?)P�Vۖ��!窋B�o��Z��|~2�J�������"�I~gc��).�"V2U��� ��]��	�ת�ۿ�L�;{&�-h��qKj�A}G[�l�@�9s���@�~�;Ж�{ؼ����Z�A�����0��I�dPc?�AY��k?Q$7�å�2�e�6�
�k��*������)B�J�նf˞u�]0��(�Am��Zr�>߮5h��(�d%]�	KIx��H�~p����J�	�N�*Y����RO��XA!�oR�I����v���ψ�+��Y�m5U�0�K�w!m���3�	���
.��#�0��{5����uTN�O�T�e�Q�0�G9��ߏWG�{V���~�*�he��$a���a��Y��*l�x�Ӊ {Np?]׋s��Tę���I��^��ȥ�׵I(��q���BAR��y��ޖ�����MK�9��2)��M��xZAdc��¡� }_{1�+Ќ�V}��RJ��և������P���C:?�y���Zb��/�m4�d�*�[|�7��{眸��9�Ě�&�')N	Ǩ}��1蔶��T}���"c��eo����P
�t�Wd�D@�� d�J����.7Y�8)?:P.����)��������mvE#:�9���Ni=8�A��y���I&���(I1�d����Lf��I��S�U�� �K�hɱuTC�c��w� "Ծ�D�>f���Z�޹