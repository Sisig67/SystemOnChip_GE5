��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%���J�(J�y0��xy?019[�9I�\f�M�����h�<�}'�#�-|���w�H� ���[8����q�JFZgI��C���5v����5�-�Z"�ec��p&ñ�O��ڄ����|!?��XI0���j�>/�S���Xf[cM _����u�b�B[�t�tJ��qI�`�߼*��8�=�|Ѱ`E'v�n���OcG[4ę��Uf�T�71K~D+��*>��) n��W,��L!	����k��p��e�q�͍y�@'
�y8�D}�����黡�$�\|��42Q������j��q�n����	�Yyf0.x\U��?�ά>����}82>|P���l@�6�-�ԨA��4��bA'$�n�zm6	˰��l��`	A�� %�o�ݐ�Do%�	!�.gŶ��J�)�$�#?@X�[#�$r��*R���ĭ.P!y���袃��}��EG YX���ơ��\c (���!�d�a��#�Z�g�����ĵ��8���%���n[���'5n�w��+�v`\lu�pSHr����W9#�r�M�_�F��<��`_
V�5��!Eѯ���\���#�T�y?HY��!Y�EY9F�v�tc
����������?�ܒu���>�O8:�x]{|�Oު
,��IW��\�IzߺS�>���.��P3��d|��&Κ䠜�ЭE�|���h7q�V�HkX���*��/��^��&�R���+_4٭�ѾT�1W2��NM׏7��/Ъ�B�go!�sݣ���'q`��X���u�ކ��;i`�-��T��J�D����G
-�6Y��9x�/D0v�S_�ܣA�heB�x�6-Ȉ[��>U��7����_V���d=U� e������'���0U 
 r=.@�,'�eȞ��G�u�m+6�lh��/�k��7��_XX���D�,`�e�m/�2Rw�Յ��x�Ή�(3� �O�&+���ж���:���^���I�&d�����Op,wn� �fQ4�ޢ4�뿽{x��l�E���1��,�/I��/8�����b���Dg�D!̭9 _h����taK�d8#U+���|��qC�k�!��9"��aJ�����V�܃�N���#I}��m�4l*�)'������p�%nq����wڣ
#�?�z�����09qç,}譇{[�ԁ�oM3�,9�AFg��w�]p�>��l��t<�q�蝛���vrF9I�S].���p�$��i�;&Ke?p���}�@H�A��9|��2~܏�[����e�.؞V�m��*l+Ce4�Z�8����s�p�*ȽCus���]oI�	hi!�z��|�{�7ǳ�I�1�_ Gw��f�o;��������W�/O-JĀ� ⻣���ϛ��5�x�PZ�2I]�l���+�RG�k�����c�8�2)�mzC�{a���
���j�\Ҩ�w2nfki�����*�qŠC���Պ��k%-�ӑ��F���9��8kc�Ƙ��*��|.g�G꛳�?+K�7J��;�&k�������}�C��OĹ�����>�F�!�M�{���l��HXX�p3�R�׎�	�Pk��h{����\}��l��`�+�� ](�5�8��_��C�����L������~(իԭ��"��N�4�P�jp-�g�$K��A,�Lڃ���eu�&tBD��~7�B�(�z���)�Q��">BH#@��N����L[-��;`[��fhJ�K2�Ֆ�%z��.sgC�q:��HŎXh����2R�C��Z�	#Y�$G��.�72F��5�b~��u�s����`W.2A�!�;Vڰ�B3WP���^whd���i�2�v��W2��H����CB�G���n'b/�&�䀻@��C�Z�Y�YiJvA&(�������"�+t�<w������d~�Ta�a��v|���9��ڦuSn@�gF�tɜ�0e�}=����£ϱ8i�u<��ҵ���p:�1Q��`��L�^�����WO�	<�E�������[\�zt�gH�@�]����\�Ұa����9x.�ȥ+?* '�Ȗn���@�d��{����qWvK��w�]��mok��T6_@���t\yl}�VR��fL�=u��W�x�z�NO@a-CE���<Əz�j���Z2|�6���ΆB�k]�M&�	Ih�l�1���#��������͢�<�Gi@�͐��p:.Q~{
�XP\.7vp�:%�5���2���R��{��!>J��'�hƘ���|+Mj��Y�
}aɟ[.�}
�I��j4��_ѷ���>�C�w��:=����������sd�uUV`��i�
��R[���.�i�������t��p�-�MO:����`�͎��?����A��}_N��m�S"�r�8 FH�-ku����H�:���=�4�ݝ�G*��J�DQ��L[
4��ƽ�L���)۵���s[ \��#(+{)�T��q��+��CDx`\���!^F.F��Ҋ�U/����ƙ7�*6�e}���E��A��_7��  x�_�U��ؚ�Q�����ѫ��ZS$����9���nM$^�!~�)H����Zw�$c��y�KS$���-]*
}ƴ���>љ�k�b^f.q�
�k�gg?�ؐ���GS��
��L)��s� ���j��#
�_2����P�b�����+!�P^��Vԥ !
�w	��^��[�]�$�5�Veޤ��O�{�_�N�W��3����X��,�^k�Q-�n~{;�#�Z���MM
����� �8��b$�����'
��H��	ȣ��:a�O���W�`/ʽę������V� 
kQ�UGV ��P�9�� j�����,O�ff�a�l�1��������_D
�����$Z�3V��{'JvΊ�k>�2���j�&Cr,れ�=�L�{�m���U�ƧH2�qDH����\K���U�c^�����c���K�Wc��]�4�4��zD3X��%�Yy*���*�
 �x����4��Mh+AzⳭ�� 1gj���:����ݛ��������J��<�K�ǅ�vʎ�b �`���ÍW�t[��C��{��QY}r��Pf�c~�$��02��F��������2]��(�B�wD�󨺹�qb�Ŵs#�M�V��te�5�3�4S2�0��j�*�|������4gk��`�Vt�!��ViYg��\b�@�[f�
`qQq����&��<�RBhK0���ݧ��cj69�	(��Ts�����Zf% �{;���1�j��5�]�h�4V|��2�l m:#��Ƣ_fN�!��4Bx�%�J�WbOJz��T��\�R��o/yj!���>"�!PJ�v���	��>��`�.�a�`�Y,׫N���b�Ŗʴ��<�k߁��w�t$�n��8�@�*���l���=��T�Q����y(H�I�O�E��tO�|Cz)��P�S�3Kh�z��EF���t�@�uf�S�]֒%���G:�g�^�������~�{˲�q�<���Yg8+i��W�:���#�U��j�n:��vt���Sj#���S �Tۄ�d�F2��A�ha9?���w�$�L!�}��0���ڤ�������=�d� a� ��y�}0�1�B`��r�V��Wm��g,Щ\�UcD�MܧqS�TU�n���̇���2"�'Կ�3-k�)�~������QU3~p���Ph1�*�����N�6��N>���y~��H0�*y�Y������#�J����%���f�[����a��U��1���f����7�#v��n���V'��o�_���Fm��:��k�I��	��]wxy��0*L�X�����Kf��f?�T�Ɋ�C��K�	^_�5e�bC����_��:@�O�bl��v�Z�Jt�CH��[�X+h>�7���u&&O�P<o9�O�T#(�y^����p���e�(����D�Am]K_v(N(�d/״����1a)U�{��i7g�;F^�3�EQa)�#}�Ab��b�a�u���s�s����ɖ]�F�g���e�y����{]/�އ�m�G�L��2���S����y��?�4��6@ˢz�@�2�ae�@�"��sʫ0��,VO����n2�b�qB�:K�/�֛����9���G?G�W�Էwߊ���i�k�ª���Yin�WB��C&f^5����lt�y������оBZ�^���\��g.Z�a�vȫ"��|��2��_��S�A(�c{�Ľ���A�c�x-P
<k������)�k�v�6�B�>��&�c2���k�૘,s���\1�F����R̻�f1a͋V��8��V�~Iꦙ�C�Ƶ�:Y���5���;�0T�QS;��1K��v�ua��=���Mx4��0��d��!��k �X�FMz�?�������: LVB�TJ�<��b�ۺ(�5�C�`+|q��b���a���u���U'�8Ŝ��u	�ˠt�g_��e�c��F6+ᦔw�(y��uÇDu�4��pY�b̽��Uu��s�8o��Cc2�|i��������r�ʔ^�� �q���#K��A�q���K�2����z����
��I���"i�|Z�n<���]q�n8��^*��_H�h;�޷�س��x�vX�~�ï;d�9��=�n��ʏ��O����t�T;u�cKri����&���~���G�#ѭ]s8��˞\��k��}�`��(�s��&�f��0�d"� ,~�Հ4���7sW�B�u?sm�M�$,Z7̞i5�6*�ʶUp�-">I&&��E��Qd�,��e�7�xeX�v���r����U��|q�<K3>|��g�kϼ]>x���N���֝gm�-;�̨�M�3YH��ϕ��������6E)�R�,_l��$�#_dj+ǗE��mKPO��8Ʌ���ht�u1�yN�僧W��87>;9o�]x�0L�|,J��)�1�u�Kҷ|~�L���