��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_��՛	�D
��أ�76ϋ)b�%A��չ���������U��W|���:;�@��V����,;��5�������ʊ̗�Y���ÍA5O�K�G�R�a��lu��ZGo�yױ�W4U8a�ے&��[eQ��
,+
 �5`im^�����;>�TȎ�i$D�� X�'�ȫ������b���9vPq��\C�z���X93��^������,��	Qi�HE���p���3CE�/K�:j'����#J+"'������R���NR�������a$�ʂs9��LD��,�b������0]�x�Z���3TKv/�(��W��pN�X�^*���*8��l�h�����R��:�ƈ����/�`��{ٻïXQ�>	\�"��ɚ\6 �ex�@KNc�M�K��[��s8�h��_4�����3V��P(s���=�LL��6b���H�_K���$��Zٻ��֪W|��m�#�2��>8>�PƂ�m^u 'Cn�����84l�'��c���:��D}��"�wMA�x^Zz����V�����~�,��xDpp)������]h�J���/��L/f`����(�8V�ʰ����(�uc�Lh0��R�M�p�&T*N(E�Y�U��\�[T��8��!�>�f�_�1)�@)�|�d�(+Q���j����{ñs���;\E���cQ��WV�=�&���mF�N�[�P�o2V��X2�D,��m����ku"�ϑ(����X�s����B����s��)R�b�NB��h�R\e=:��&��ZW���F߄�E�(F�+��"�mO�.6�s�|��*}��!�ޝd��Q��n\]���~֩Pp����90�!�a��+S����&#נ��BE�!�[�K�+MC�gW�t���§j�Z����:�v�������(�q��1 �s'*�X=[p !%��sr�X]����'�qj�]w�ň˚{�mA�%5��K��0NK��@�> ;.�Xx���/�ص[�3� i�m�*�6p4"�X�Zs�6�fv��θ"�5��(�S��)$�ј'%?b�P5#�j۷�B>ٕ½^�7ݵ�����;^��Ou�(�j_���EˊG���̎Lgn78wA�+p]D��{�]�m�ݙ뢐|N"�6Rd�t�r�S��W̚�7	��U��q�ܻ��|�z��l謮vb�W�; �5�>k��+���؂��*�%�nR�B�r�m�����.���.|���4yǏ7��V��d��m'�����s�.(��'���U�N4����~�/�����P-w�fX�ަ\.!N��!��<6A���"��B��C�4N��B��Dq���:�@�*��� ����ك�thY��)�*jˎ+L����xuR�O����e��ٳ�i��	 �R`�qŏ.|�P=��L$����@q�"�4�u��X_��)*���/�T·��q	x'>��=$x��B$Y������}��#�G��_o~�;x����FT�+Rݠvj�P	,a���L�v�9��B���:�`0���;J����*Cj�*�9=�@�� �I��j� m��7�|ٵh��*�T�y{}	����8� 	T(;��BH�
�H��w���0Ad%1��E�l&xvJ�	̖����FY5����٫=0�[�H����=����8��\�*��Ə�@���RtE��O��H쭊/�ѻ6��U��s����c�_놙����ET�%��(�#�m2w_@��8j� �� L߸�(d���z��z��"�؎�%���8������`ݝT��6�tc�v��g��2f��`�v���L�$a��v�%=������LT�*��r�w#�3�~����X* 1�Ʒ�{�0����<Y�s�qH@i�Pv�6����o��� Ǡ�&n�2�!��.������Wr�:�t���\l�V�+xb�"Fnt�����է�-��ܕrE��E�W�
�7�i�*{�b!Tb
��%�ob���c`$�2� �U�G���'��a$Ax�hܺMo@�Q���v���4�(�Z��� ^+M����{��S�Y ���.`QpX�E�Vu?�Iv�*�y��0%�7��mT�$8����c 5�,���JMuZf�s16���j�ڌm�?>JZ�n�Aj�n����D��X>�����}��H�^�}�<ۤP|	��&|���.�	e����E�����ז#�T"�����ՕDt�;�΁�G�X#�������<	���(�ㇴ��_���fs�:w��{�����т�Zf�:��<��*�����Q��TS�ꄤRq�a�Y.�3u���f�&eӓ1����ኹU�p�d���77\����[���9E+�0q���#�_Lf%�O3�ǱQ8���DXj�2���=�N{��+�5�׳+q�1�� �d�\u���eB�a����x�T��m���Rn~_Û�x���B����VI;���Uc��X>���6'��ћ#T�t�R)��~+���Fjq���{&�ɾ
@���g�d�)3�GRR�K1����9��ޟ�
}K���P [��^4 �N`�㧓��W�\��^��Y��Q�De>dO�P<�<Ӈ@<�kt��D������։�b/ϸ<��T�9�PHi����J��ȯ�ٿ.�E�(˄7�O?��/m(0�m�28u��/��Fٓ��Q�tħ�g>>��Gm6	j�aP��.��&��gE�+�s�TM��H�����	�ڔÊY'e`�j:
;���;��0��f����� D�GK�L�90@�-��b���/#aKk�~�����ucڏ�Ⱦ��xk[�$.��@d1
��s��^���uzT�#�(�i����c�Q)E��د*��� �^�S�薍�I�vYƢ7?���(ԃ��ҊIq�!S^i�P!��*�
6��`��Y\�:�vI��JBSA�}rN�Ϋ�pL��}ܢ���\�%
h��6�<�N��֩���B���@�vСl\R�RWR�dm��	�8l����W���T�=�q��f�!*�9�8 _�� �����lpF5_>�i��v;p��83R=*�Iw�˥B�I��O���q���]@�L�Һ�h�e����d�w�q��S����r����Ƣ6m:Q�� ;���H�@y�B���Be�*�T�	���!��l�M����`!���_ZA;�_&�V�(Iϟ��Yn�x�>��Z�Adc��r��[��n��d�$���nkv�ɍ�|w"M(M��-%Z�n���Ų��I�lRW��!2q����}{`�4������0�7D"�&XF�? ����֚\x{?��H��%�͒�?��rcQ�K�vU��&-��śh>4U�t�)��Ϟ}�
�4OKc(��E[��=�NХ�sy��Y"C����&�&_�l�Rك��`���ݬHm{WE鈔���C�Hp���&1x�`�G�d-�>���Ғ�ҙܡ�Z�9'Q:l�D~@ 9ts�Ȏ�d�e�����	��+�-�Y����U�.X&�BEa�tmî�]��Y�3Z�l�G'��m/*��,� �����5t��ղ��%+�,�	ĸ��L���K��e7"/C�5���et ��7�Ĭ�G�ulĦ
����eFBǝ 
������C�����	0>fz0�Rm���7�'�u�LX�mB��\ r綹�g�I+�1Z�w���Q�� �S��:�<�	)=��}+!��M�(x���*�=k�u��m�I5r�+�n=3���څ-xO�9w�s�| P`!��{?	;�"��eF�9Due���W2+]��O�!���R`�c� ���O� Q٨�h��o_ى�,�N=�5:���J[�>�S��X�������M�tL�=�� h�i��V�3p��>����z��Uˤ����o�t��-��!,�'+��8�U>A@^$��&�#g���Ej�9�EG�8��Κ��*gv���`���D
/�ˤ^�s}�^#j�Q��9��LQ��:p����©�tI��a�᭡��y���g B�x0�a���z=�[� �|a�&
���q�r��P�'G����-��LU�������-O�kl.ƱCi[���~74'�8���Gl���Z���"��yA�,V��0x^�G�"Q��B�2�=o���VF�>p^`{�l̔�1AʡA�z�V%"����|� ҏ�=�3�i�z1�S����,*�5�V}�����xl(~�<~�u��WW�i=c�����Z<����!T�=+�ݻ�.���� ���l��w����g�-�h눏k�/S73�-����h�t��c����,�P_��nx�/[8������ǐH��]���x4K`��(�*��nstB*��+<�=f�m���3�j����uE&K<C�?6%�ٛ��k�2�B�`SG;m�'\A��b�Y[Sy$���l����]�=S��>�*PzOiM���!���� s�p�n�V?o�¹�GW� �H�S���{����&��e��V�������@iY9ȼb������*~/�R��ll�g���2�y��iMWe:�
1���V��8�ަ+��QM�҉MK��d���r����<��#}t+��3n|p�[�N�@#I�V<-�-����2ũP��Q����r;bl�un�3�����k�7V�Hs����yz��+�]�=m͆�ϱ�ZL_�}m~Rk�-CSgפL춓�n�b�BA2W��J��!R*�Ļߨ��o�����u�(�(��� 	��Ԃϭ{d\�ZS�)�+�S��{��� �Z<�\�O]a�D�N����O:	{��A�ҍ����C�Ÿ�R�'�u��~}�P�,����5N�Cc}hf�\4lc��P�J���&�t��W)�&�?4�l��7+Ԋ����Ez���{L�pL�u[������U0�+�ں/�-�3HT�:��	-��ņj��J�	�̿>�)q~��H��������/�NE�dmQ� ��,�����춫����?��C�0f�����U"q��p]Ep�ڦ�b�!��0�1�c335	1�-\�S��[��%�VR������B�M�H�N7�Z)���k���4 �yV:0�Wό6�Be���[���� ������G�@�V5R�7����}Z��F�ʅ;�(���΀g�`����>� A�	9�%'팑!��r^HRy��0o~TN�<�ߴ��)7j�<�r1^4+� �(Q�<r���:���yȢ�:Rz��<��~M��la�8Ao���A}ވO�*��|wK<6{O�~���B��k�pK�E��}~Sν�l��х�����j�!\�_�X���V/��1�z9<��a���p�p��1&�.9DPt*��'ӫ�9�ᨐ8�۴�\S�ǒ���,&�r�]Ky�}P�<3C[Ԟ�5fV/����}��n�Y��6�ќSi����J�ʏ9��#�V��$�e����l�u}[�%�������%��shR
�;%0�%����f��є#O0��A%C���G�Tn��n��₃V�	ӥ-�X1��WX�����7n��I��,|�M�B^�;!w�BA�dz��0}�]�jwΐ=�l�ٴ�0C�-�5o+�|E��i6|}���sѷ}��N�H�҇���c�ܜ�ñ{/Sd�]t㬂�H'Igg�̜�<7�&�ѝ�"��!7ք���[A)@n���aZ�hڑ.;�Y|~��}eG�:����5q�)��d�%Ѵϵ�&�S�C��ĺ�F�J���(��Q�/<�T���P9����a9[2�ni�~uܝ1/� �Ό�l��٦U,\J��C�Wf��ㅱ�e��jۨ��#��y�d|��Y�=�nm�q�1wty��P���x�A��1�b>���]��2u��y�1��R5b�)��r����5y%�Q=�	�C�25$$m�kbr$|�*���Mf�Nt�'��N#ʁ��y� Ϊn��VQ��/V���)�bb��Ьb�i�B��Z����+�����Ō����K��Q��]H4Q�=E�2P��Vޫ�5c��6f�.���r�l�t4�n�awM��(X7�.=���)_ˌ��3Q�H�/i�P�
L�aTw��R%D��~.B}� ���к=pv��"��ϻe��Emh蘰F���3�®�q��g7 Z�~���� �6B�{���8��C1�Q��x�����򛣺=�����]$�wv5{Gw�5�zh]�x9��z��S�n�-����s��@�L�n!��MM��!:W�J�s��!hb��[���e�*��S�];���]v+'p?�?K�yCNC�u�*�<��w�b�ϳ�#�E!��q�$3R����8\CIƶ�u���y_t�a��L��@t�(�I�����<�*T�����MJ{� ���Kʃ�4E��AO����J���q}e�w�Zc��P��Z�4��Ԭ�=)4.���d�믖�m��"/��e��XD���WS�_�dN��Ԛ���9	���tg/�r�n�eAV�,���.����8.�d�#��Be�?m�_.��βCa����ʹ�	���X)=#.L��<�e�3�����Nt�o�Cg-�O٫q0��`aB�B[z��+x�7�i����$�"���_��܁�lYB�vq�\�5��^r��O���'��tN
,�Av.Y���w��ePO��O+u�rгLӆ�f���1����L[>!��!V0�$�?���y�6�I}Z@LӬ�]��#�S)�(�o.����`-��Kc�
VU?.��/�fm���k�Ӟؼ"�	.�/n`Sb��|��13��1�^�֗ͭ�l.to#=��kBW/փҤ6�뵞����i��F-$�lpF����ҕ��Yq�羗	���7Tb�4�7�Y	�ʿ>�Q����Tn9�
L-<�n��"�S5�I�Ŗ�؞�`��'�U
�Ƣ7|���2��o|�AI�uͺ�1�I�������2�I�,7QYR`��w�x-���B���3�`M�8rߩ}�v��'��s�]����,�Ԝ��LW��P�4ġ��r�"�33�X���uЯɾ4$<��0�ih�-���p�5'���F��L���+�Vj��Jݷ�.p�WZgN������g�e�^�ٚ���l�~�L��[;��[$�fY�Kb1�WT���cm�FuE��\D�p��ݳ���,����O�C��btҟa{�.B�K�p��j�9[;[�i�I�~��N~����d�{cX�~��������h�.�2c��s�84�T�.���<���x!���A�#�k�B�`��?�1R3��V0�Ë�ns�G^�T������4��� �:r����1�6���޽%��Ћ��(_#���,U✄U�=�~61v-o�<O�$.W��i5SMR�ؔ������覲�.�-�5DCךw�p��m���{��z�G�";�����xq�y|ۋ�x{ح(yF�R\�.���b���b��<�O�,���OD�:���;��D��KC���%���T�ų�}�Vz`�J��)�;�~���P72V���[�>��o�c��'Ӥ�4�B���K;b͓��0҉��C���2��g���w_����`c޷m0���~s�I+,	��$�I���<�@�k{� �C���D���.���MB���1��ܮ�}��u�p �ɞ����Ň>����Λg�k��!���­�T:i�d���Œ=f��M�ҩf��>5���|�hdf��F�!l{n��X"oD �*�t��d(��Z����#���e:}1�}���l��������?H<>Ho�]��FQ���
����L���U�4\xh5�B.�q�cLq��n��^Ք%��I��z�Y��::}�m�u�C�b�;��{�4-�*i槹�G��EB!84�蒻��I�5^^mm6,Kc�G��:_��-%����&��sNw;�Py �g��mx�������M�F�3I��4)�gZ�[�6a��'�o�X���4�����ط6#A���%d#��W�֐�\ZìB�%����-ﻷ���Q�
���s��:�������;,�5���bY}�7s=�×��u۞¯��X�Q�ݸ�1Ԡ;<�B�"ꆾ��(EK��H	��z���l�E�\�ؕχ����f���r�ٗo� �u�<���>��q �J�p����(����"���@.�yo��ϊ�~�(��f����e�.�%�zRdǟ��Α���2�&����s i�$�!ˮ-���pp�&\)O>'l7�o��M��'Z��Z�6�s>��|.��t~*A�\��ڐV
�X�,�._ɒ���aGG��g:�iIErX�u��ѬHJCbS$���W�n��],��.J0�0�E�����dF5M��NA9E��>r��L\T~9)vlE"��޶V�c�����m�	��᪘�/��f
Ȍl?׏������	b���עX�6�ص��&��Z�|[��֦͆��//u�<��I���*ݳQM<��!�n�������x1z���<�F�1�zI��+M:�����T��/��`Re�/=t��u�B`��nd*��z�-ڻۖ�fp&|������F�ڿe�����ʀs�~~ �x��4� fk���RɛS�Z8�T�ǪY���m������^���M ?��n8��M���A^Md����u��1�)�N،�+�kO�0�+� o ^W(�m��=B6��7�5O!�,i"�3�d����S�mNl�rZ��6�w�xTBEۉ�������%� ���������V�#-���!5V3�|�l[��b�h��\�'���)�@�zҚ��Wq�"�6ɕa!�:l�@o���B��lY��������oPv�w�=ޛ:�RI��5�	�E�6�E�?'�%�',U�E�>�'#dr�,HD��֤wI���Ź�у�,� d��R��<f�+TS熱x4	�@�"(��&�����O������}����ӄ,<���@��d���.b��epic�Y�b�_q��$��.r�`���DH&_�x׎Qh�Qu���"�VI\��0	�yN��Q�"�#L��ȿ�2��"oq\T9q\%�R�0oH�-�Ը���K��X�ǩ�����(�)O�l��l=�����M��u@���F �&�x*^R�Yföc��H����;�����䃷P?^�kl��n1}����鄊�3��1!D�-i9}P�pr�� �y�%=ɉ��c�[�5����E0e`��׹$ 8���j�oL�E8�n�͘ac�h�P�=^�S2�20;�}/A
����]����U��Z����i�@�&��^�*��+T��"4�˞��L�S
�f߳�m�I!���U���aM-+�� �BAn)�a�E�$HU��Ռ�<P��:��^u�IG8{�А��}-6	��s*�'�D.w�w���`� �	�&i^�S6h�3:=V[=�!�u��MJ���'��x�̞Z�������5���U��/{��n�zA��̂E6�`n�	�x�}�����g;�6_���/y@��X�$���j�h�3���m�~��U��Ʊ�����D��(g��a=�N����3_��0O�8ݽ���H�N�W1 L]�>g0[yN?%ɰ�1A*kS,���ivG��fF�:� M��@�hWΨu�P�9Y� ���e]4�`Uӵ(1Ȟ�h�0vEu��`��X���)0�^��7��<5�S�-���I �C _��8�)����x�`c���K�F��/e�Gb?��w0<���U=�f��`~ ����EP�<�p��x�?Jv�_�Qd�A{ꍜڮ�_ս�d��%"�E<�҄��6��2!��@M���M!����uf 3�`#��g��$O,�SGػ��ی�Xk��넘Lg����q8���:%��PR��ih^ث~�.g��`�6%;���:�6��(���j��􂕜}M��ŮS-���eW߬ �V�Q�]��f�}/)�0(��Pk�A�ǒ3��^��E�:U7KFu%�'f�cAA3��!,�U�	+sǮ:Z�V�dc�΢ \YP���
�}\�tH�h�,�!E�Vi1�ޠ��DS�����ET�fZYH�+֐�9��ҏ(����t���?"��9j4����e$�Lt�*Rpl��+��-���~�G�T.����G�{�o�G�����̓<r��<���v��0��r�B���}7��I���
�>��&�t��9�b�4�,';5qH�ˑ�GxNy�V����3ӼL[�߭�D4�R�_R�L�M��֐��.�rF��A��izϗRz�r8?�o��JMN����"�����ꒃ�~㵅��:=S��()�hT�:�r;0�#��0���=��:-��u8�}-����sh���csڌ�a�$N�����e���#��ؓ��#%��
}{4�y��ۅ ��4M2���s�4�V�;����t��B��r�~��{��?���u���.�����'ó/��I���3��E�b�@-���c�Z=��4e6V
�:j�J� ���ߒsx;xG!4�h�+D&�,��x��o�Ր�º��;MF�$8�n����'/R����(��Ӣ^t�E+SlX������mnߦ��Pl��I��k��/�ڮ[&]�]ZV�q�ѯ�`��4�)��1p7Y�A���c8�:�Umo�xC�N���9��t�����Jh�	Wob=hˏ�$�w��޼�4��b�#���	�����a})m�>)A��m��ڗ�a�:m��`���5���ދ��2��S�.�RH��)��~��Y�h5h�F����y���M;$��|,2.Q�xРy���,��}���̉Vd�	�i�
��t[%N,a�yAK�"���]�՘�IdT�d͟qu<��F����ě>ݩJ�	_}yn��{�����ݍ��0�S����^am��N�x�E��"��,��ꋪYS_Ȫ��E�Y����3�ҷc� ���˂�js��<h�j�������!��P(�C.>|�p�#��FH����{	|��n�u�1�2���#6�Z%��c�.Z�F�٤���_/��S܋(�@�c���$����kB�4�e-��[�zs����c�zHd�}�{<��,@���|��4n��"[(��1��<��Wqn-T�ܫ)�/P�[�u,����jC�ۓM�Î�bP�M�g��~��nGK�G|��**ߓT��W\g����H�p6Rz�N��h߸�FủJ|�泃GtM�����Y�q4���}
c�
��Z��Z
� 4 ��Q�H���RN��H��=%8�l>~sJΩ��(���@�$��C2܇��;M�� %{��Z蔶U�l�-ѵ�u" U����%!g��7������s� i'T�������S�жC�+��'���Y6��l��t�)R��A�Ƙ(i�c܉c�h!�o�h0���5mא%�E��9���_@G��I!� �V��/0;t:űґr�>3�H�6ǯ��?zT�Բ�����̵�T �ԓm$õ�T��W�AJKk�^Gh��gmɾ.8o�b�P�42��|=��t�)�r��`����eO��0��3�#���f?�$�r�<yu�'3+����gM�� ��Q�i�b��z�Z��7�m�:�;�}���༭�;s���5"��T��%j�ՌJ1�|#�N��n�'�\7-y�J�V�_k}-O�s��B�>�o��r�|>�9D��j�ao��-׀j����q��.��$�X��rI�F~��j��P��Ovn��hD�2�
�C_M��Ԩ9�_�E�=�h٦�[�36��N��v�s���n�6���=����,�S�<-���;J��<o�>�2�����f!p����`yi�X*	�e�-�����9�6��v(����~�P���T#�f���$�ڎ��Td�`���6y(���0�vE9��\b+S�����Q��eQ��Q\��l�I��ŏZ�����5�;Kl�,my�s����ՆS�tc����~����"��:�Е��"��3Ŕ��3kiզ�U������;M>�n�ls/m�W����c_g9?��|b�uOh�V��N�`\�����;��=�px��:�G��(Cm���>V��ӗ
�ș��#��2��P�/�:�'{�>��Jm���=��n�V,�$�޸B+�.�x䆳�]]��T�J�V-�0��Ű< �W��X4RA��'�9�J��.�a���F�eB��L���9�L�*롪��F� ��ޣ��CD�\�3�vn[�"���2d�i��B�H�����C�p
^=Wf��A�\���9M�F5A�>�%�.�.���?=�8 �  Q25�>��x�+-gr1OEc�c�TrN�:��TD�RP�9�'3V�i2��A=��s(�T�vx��P��Q��x���$�������x���\c��U(��9,��lh�<g��	�2�篛3�WFz��皒P5�R�a��h�TEMȕ9���]�R��x>��Q�
�^��PB���w	0Hj-a40���k��s�qƨC��wQ/f~�����Xb|�������R�?et��g~���[�_�JQ��PS�]��I ��Ch��͓Ո���d�m�2�/50RB��� u�й7��
�{\�Ǧ���$�A3߉�	�)�|�Y� N��<&;� �>~?8h�S���`�#�}p�o��	jef�i������j�Y#�������;� �9N�b�8��2���W����)|>�^��I$�y�p0�F��FrTcR��1�DSH������t ��c� bH��]��A����<C�Ɋ��q]8��`z+<�WQk-e�>ic5Z�h~�b�07Ɖasqu�I�L*�g�L��=^r"�a؞ҟi�y+��1����1fOJ���	�4i�mG ,������Y�YnGc�x_��*0i4���ZV�|����c�� �k�o��b��>�2��D�&��;���^��2�.�O�n-ʅ���|�<[�Ky~�$շ�n�M��փKv�4��`����k�U�䗋1�ڷB�*U?�Ԗ]n����yE�$��Y��>�:�Sx�֝����e��وmؚ�ۀQ�QB�̞�#Se� �m'49$�Qr�k����Xdm��Kz�����"1F��>$M@g Ԭa�� s�\��|GD����6��ڨIp���Sv�΢��
o<P�6�w*�.0�"��\�N�f���>����6+�tG:���Ԯ ������N7��3�5�m������Wz���VM5�`�3�(�qraWF����ӄ�S�^5�P���4f� i�_������x�����o^��	�S�-� K�G+��!P��4_'.������i�lp�~t�Чu�3����cpAs�*�\���3���]x���9��j�{��;r^VJ��G�[�W'E��f�#�_m��΅���m?wRJ�xH⎀������'�(������_��P�}�i�Xr��6��:���܃ ���c #�^��w}�b���#���U�-���-X�I=�x��Z#x������Ʈ�e��2i�#Ƨ�Mc�D�i����Gz1���Ab�*���Т�*g`*�Eo�e�W����=1��y��Mj�}qYʱ��I����㑮>o��'pٕZb�[A>eY4l�R|��,���ot�]���`i�mV��g���c�J��Bdd]��#�_���]�=)��M����F���%�6�-UoG�� a��-PǼ�ܯll�x�@��A��_i�����ڍ�e��U�c�-,{8�s�XQ>F,݂�;"`��۰���4U�f������^�g�=*��C���!`���2.(���M|oԠ��@҄�D��)��l�am�\>�zSף�挸��keJ�>���Z�rn$��͡^M�J��ٛ��ihJc��~E�u��8�(�V���5�u�(����#҆�`�<��8ؼ(�/����C�ܚ�z �ͤ'^狜��h��+�i!V�d]��b������U�ޕ�z�4�,�r�N
3����l(|f��).W?j���X���gzg�2�=�d��ŁBt�΁p����''�jEh���*�A��� _T9bf�~��~_��	��\צ>$@MƁ��iEO����M��61|�����g��Л�L������x�������� Ŏߒ����I�b?��U�a���a���r"E����,*����mH��c|y��x�z_��.�U\��(]��GhyA����2���G��"c�Y�Mƾ�KW5u�aV�����o�%4����p����CB�f�㜑F�0䡜 _k����S"���f�j]�N@8�;��1w��K�*Z(TB��/%�>2�j.���"gL,�orgRN�I��p��|���+��#��[�-� ��Z�	��zқKR�������N����kB�!�P��tϒ�EJ��,����4����p4�F��O���Ukc���'�;��?&���oF�g?l�9l�$�|aS>־�$�@�j�-�<@&�S��X0nZl�p��P�b��8JG~�add��أ��|�:x6����S��
�O��(��I[=��d�q�S /G/A��:�R��V�3�ձ�U"��F���:!9�b��֨صЪ�n�v�V㒜HCHK��%��Vu���Z�ߎ�R�'��n�&���� 0���%ʜ6��V-H�oh���׉o� N"��l��y��*�<�������-+D"r��ޛP!U^�E5@��9&P)�����|��s%:R~���{<fΪs��ր	��Ϝ���e�o����knNO �ƙ�����"�
�J����,u�S���P	~y4x�Cg��=��c�^]�\֯L���9A�	��ؙ�)�塩��<�_;$���R�C"+Kh����`o�b�4�J��/�3h9.��f�f3�������E��qGjv���Iĩ�<�7���4wjN��C/� ށ��]�1�����LW:�
����ʍF>���Pm�7�p�8C�����O�t�	n�"����P
��x�Wo屹L�.��G���¦.'������R�u3�)Y_I�v��Zԅ�gf�D �?h^���8j�5�s�k�#;��iAfw����bK8]�J��|zHZ`�Ktn�	r��M�C�`�²K�0�\�0���  5�j�r�f$G��	��C[�o6a��2 d�Db�t���ga$����'3�4R��\�t�p����&��-��|ܾ�D	�?t���sE_c��Pa�B���]˧b���{BѶ*�d������<�A2����uMb�;q!FF�H��f�T���JH�8)����4��0<�yWV�R4w샏��*S99d��&X��\�q���ݚȠ@�P�&X�Poo�g��Լ��ϱT��@��)��@�/(�L�ѡ΢�V7�n	��5�Bɗ�G��������/{0Nf�S\`�d{6���؇��n�3�FUs�nF��Т������#����<D+ע�{��O	���|��Z��.x�cH�b������*��j�]��c�:���u{�S���rM�)yy0���r��$�iu���W��v	>��R���:"���;q���bb��đL�W�Ïa��J]G�S�.��,&shrC�0X��;�������Ǟ��{IbCM�@'�����撿���t%�hZ�A����w�%�[l�'����US8-�&Q��P����byz����~f8�5@v�����L�l�R��TgN���2�ӄ+a�tу>�#�����h�G�]���2�̰��7�B���b���E���<�T��R���g%��@�����EX�^����Z�w\VaH�]�� ;U���`^6u������&n��������%y='@�dd6uM!��n�����4��-����d���KFe�]TY�����& հ������&_ʅ6�2��'��{(W�L6�q����ە�/Y�|��jx��dSlI�T;Q>wƸ7�&�.i|Usc���֒�GK���#Gw��^�t��Z��{'ݢ�QvX�bтWI�j�3���<�]�eiS�l�(���� �]��+(�U�_O'B*eԘV|<�-�|iPu�#�vm�)Ym��/�ޒ��쪔��1�n��&8u~�����^��ԛ�Q!�3�_DJm�B1� TY~O�L�x��J��#�"�K#�N����+8�)�Y_��4aa1�� �N���\X,Z�����QJ�~���y� =���� ��=�Pr�>�8�̺/t����`���<G�@��h1��*��NR�H�x6��4�&�>�~��"��';��]V��xWꖋs�S��,T�������:ھT-p9���R���1�3�>$X��=k_]����|W��|���_@@����e�s' ��4*3�+5�<��m��n�T[���b\B,�>�=�{��J&�l@{�A{!G	��ޑ�������U^��C9Y��IR�i��I�i�h�#��H��ЙI-"��OOă�ql΃Ч�n6���W�Ԙ4-Vq��J���+���Ň]͙�z��ݜ81���ӄ�c���\	1���;=k�Ffo0G��# /�ʖ�א� ۩�t�ӞކfkFx��UX�����+�#y��7�M7#�њ�����=���4%&v�w@Z��S`P7�\�X-�Ow	�zd�\����
��j�^�����A��x� �&��pb��V�5�{��k`+.4V���ɁMjx��=��ilBK�Ȏ���)$e��ۚ7�Pwؾ�I"�9�E��6*ǝK �l�`8�`�Y(�:��~��L�͇��A8yݠ�����8Va'�J5H]�������U��y��\}�����~gU-�>	Ft����# ':�_n��:͔�V�d����[�O<F\����k39j�l-���_��,�"����~R��5�H�x�ح\��
���o�y�9��jM 	E���ek�8�(�*���i$XY?��H��F4r�ժV�W�> -���I�J�['��!@2yD~��*>������t�K�N^�Eg�fћ<h,H����r�m���"����͒���I�'��=�ΛBdLU)*[!�ˤ�]��q �&��t\[>�Mv�@��œ�{�Ez-�@ߵ��v��d�E׸���>č�gQ��8ר9�+\Ao�Bu
b�G�ԕ�* �]�p�u"�aa0���d�r�+ie��Y���E�Ƭi8H	8M�2/yF�ع�����<��Nnl�QY�Z�U��r����˷e����*�Ck��=u��)tN�eU��@� ����a4��s�n��!�%��e) �Z
��4��|��hal=��s��X� ��c�ēT|s��k��5����:�h׹��8��[\o�����!�3r�H�qM����ȸ��"�*� ~����'�-���>����e���f�X|%�|�#d@��Cg0X���L�SʃßVϺ��)�E�-���U7z�(�.���*}AQ#Ut��o�
T�6�b�����ym�c�'�	>�^e�)C��ZgtЦ�h*}zt�h��Z�}F�v�p�X	
�9���W�m�k�����K�V盝��[�cY����Il�lt��=��ʕ�(�XxZ-�fO�1DT׽�����r�v{Ri40�4o��W4���OZ�	������Rs�+�d�6�י�#(�N����lr����NB��:W�[=1�s�����}���i�"}�刭�� �K����	�GFjs',L��Bw���-�l���K�LD�T�Y1��p�}mJ���[Hq���f�_@>wH	ڇ�Bh�bo+M�����мj<���ur��py*�@Ĩ<��t�>_t�ݎq��76�p��#������S�Þ�a����6������[����,�P)�߄��|��h�3�A�<��������2i��.���lp����пD�"��̓�h��'���q"�"�z"C���'=�&<�.O�{0q7gJخ?�K�$����Ec|���\	�uͼ0O!�>`��K�PD��������O5���ժ�W���J�������ls�"^9t���yhT�.*����3���Wv�l�� ����el�i�.�7�n*v�x�Ne��ZH����I�N\]ˏuU�@$B�17��wo���*�B��L���2(O�ÄԷ�y^��I�?���
�d*�M��ZjM��^�o�E[-&���TdR"�?H�w9��JfoW���ˈ�`8Q�̺�Qvs:`�{��*������0m�.����������LHZ+�U���4簪퓛��W�8�%,����}�q�5c{j�_S8��X�S�TpK��L��^�6d���:���#ŦGPF��.�6y$��7{�(�]њN�AM���+����7��}#��"F�@Zgå� =�	b�FqEF\�y�/r��_�kc����:M��פF�oPЗ��΅=��3�_]�[�A֞t�q��3:��b��F�m�����^u�du>����ǖ�R��#S���F�xEFVt�u�&��n�/U +����k����ͯה|~F'�â��2�Yh��d�d6�ۭJ�rՇ��G�ؖ�Ў����=\���v�����P�����)��ɿO�X�<���q�!�0k���k��_Z�}��9v6=�2Q�sj3�%�����v$�U�����OSV�(�F�svy���;��0D�Z�K�4��l�z��]���x�����z��8�W�H��@M��-o�I_o��@����=��9�(�T�)*WX�X�N-s{(	d�	^����˸\�4�Q���su���	�A�V(,��a���?+f^m�E@���=/��r�KA�7z~��۰�.�/]�
$[?!3v�y��`��vE��Y��	���Q���U�P���tίan��%E��s ߆��$E!#5�e���G�T�=�����
����Z�Ӛ�o䗶�P-��9�n�'�[r����^wy����"�	���K�jx�a�&*_�l1MJSY"�{c����G��x|h��K��<	,�_�bo��f���������+�/���nH�aP*!�mD� �e�i�eHl����Vhue�D��|����5-]�a�{sE�=@^�-Lvڦ�!Y�@�zM�S�ĜuJ�~���70 �ҍ�|���jy�qT��i7�
 ��4���z��t��S�nj���z��=w��
�y��x���׀'��E�Bt�ed�ܤ�7�p�0�s���\fZ��Mm+5�q� �X
���4�GE����Z~<�����wfXg�8qZbslj��!��s �θGp��WM쵅�@E��W��$i�B�qv����.TS԰4y��������Քx��
G�FA��ch�K ����G�*��ڗt�m�A`J�^E�N���Q`��j7F�ګ��"��h-�Z
 ��m)�Z�9^@���H�ߒl�@�Ә%�^R�D��wb[f�E�iD�d2U�9���3���T�i?Z�ŭ�&��NNܽ�1�Z[�^]w���񚻭��JmR��G�~��`Ă �:+)�P�Q�b7�է���{���@��<�ė}(8p��;�`]��%"/ ,�0(E$e���?�$���Y��a��+���Lyت�����s��K�k��)kO�o���kq�cԫ@���;qa1�	�keR^��0���V-��4b���/~a�1l�-K�7F��<�����$w�~���x��&Ι�&�� �(�=�E�O/�1͗������	T�
���+���-����5�G�u��l��bI�����q���$�:P>�iѝn�������7�^F�5�s�0}H�ظ��f��>"�����w���[J��#�E�<�$�j_���|HN��5a��E]��`iW��W����ck��n���@T�[6Ǚ��%Q�a�5�~�@������>}P �^�^�[���,�q�j��/��NU8Z��o[4;Ua�nq"
�MI8�����������BN��6��[�Z��SIEr `�46=.�e%�]�7w��n�Rizb����sᷱDE~&K���̛:G7�L����j�44��j��ǨJ��V���Q��(v��"U#
��U���e�/N))g�
���f0���q�����t;�"�[��D�u@�R�K��PV�]y�,�e\�6W������8H���w�b�K�|NfIvY=Nk=d ƻ���ҡ�,��q<e�o-f�`u��~қ��p~߱����Aj��9i���h�+���u;Z�@�Ir�w��E����3��"9�^�"�c*�R��a������'$��-a��|����P���;V �/�[�C��-@�'}�,��U�Y�܅�ؔ���Svz�.(Q�?�ށs��._��\]Y-��kg����M3=��ڊ<ⳉ�y�h���3���T�2���O�z�<��yB���)��&LT�޻k�����#ڷ�K ؎m�gNݚ�r��\�T;h�ʗ|���'��e$�{�HN�$XSǛ�TeD������Iu����MI߹���:(q��A�k��u~�����,@�L���R��_�a�讶΍����ޙ������^��\,MX�$`�Z�ˎ�Fj"M.��_����5�kk��AUt�����{���G����x�s�:3�r�q$J-�n�a=7)eM���^�a�p�?F>n�D�^���>���>���Z`���x:Ī�t?8����q+�U� �m4��������t��ԥ����D�� �c�LҴ�YbZ�_�	ilH�s�]lvKT`|�I���۪}����ü3o�b
� ����
���2�v�~�Z>:}�<�e�S�c�GՇ�)�ð<FR���zPP�5R2�C���3�Fn�<��S"������٣�/N�VJw�Z�����)��|s�Th�}�ߴ���W�è�Gd���l5j�Ղ
��=�	^���0��6@��������8� D�C�Q��}�}�=��x<�C�_1��u/s�\{�8ڋ��O��-zi� 4x�V�Iڥ�]��U��@�xš+�$U'�-i=i��A��{��z��mSDnW��������O���}&u%X�4qn]��S!�~����l���w(�������#/фp'�����cS��ɴ�����S{��!e�/�U�ײ!&q�ܓ�����7n5����>��&�A�F}�^�aG$�=l-�m��ƕ�+�E��{>��L��B�i&v�JR��c[�p��$�O�/��)	f�M�P�y�C��H���¢Z9Cg�Q{�j��%�P`(	�>�kv���{x[V�S����L��^o��%aO1�����"7��]�?Re/n_�<j�~4�.�K����Ȏ@����?hb]D���*�C���M��
�����<t�m��w���څ�O���3���i�%<a��-J���z�I�#�����d��W��4����Nm�H�.�����\�%���ي��u+~$.M�:8�;�T�����;��DA?ufv�r,2��=W�/�	�K� �gaF���|�� ���N?>i.�h'<(�S�R���V�p��.�z��1��	�עi)�|4�B,�tG }���{\�eB^��G��!�[����Ŷq�E��T~o�	����0d�zF��#Xa�	r�Abʢ�BF�5��#���hX��z�%��@��8�U���(_JP춞��*��vP�M=�7����<��vnzߟd:�"K���TT7��5��s�Ewh�F�@�� }��H�z�5�P��e��q���i�n��N��J�����fJ�G�E}�F�$M[�j�5�a *k?�;�R����_�ޯ�2z6O��ı�ֳomp�
���C�bT[�3D�J� y�#����q ���b�>�� �,��KKy����p^�x�@��o�
������1l�<硄C��� ����P��Ѽ�X��z��D�s׊��^��y�}����2Vt���%���r�8��{=�T�wy����КƐc�*��6�o�� b 43���z����{ұօv���̀�1'�"����^#c�"$�U�/��@�C폪�N�{=�����?��	��]"�Z��B#b��5t�x3�*l���e]_������-<� 5��Jll��Kn&�J����U��n�}&.J�YlPE��������j�۫lk�p��]��6�B#�5g�
^ທ�8���຅�Ǥa�I�ȭ,]�z�f�kt����!���즔��	#�L��N'�|����X=���A��Xo �~��[fuy[H�s���_5]�D[���B#	(۟P�3�Õ�7?���m���{EG�,��ɢ
W��p�Q�~y�gW3�m��3!G�f�:�JX�Jl�QDZ(k��G*q�e_֝�#Q�100h��N���
żS�ː�Df���;���+��1&�x7݊�欝7�Z��Y��*5@A3N��!^ia$��iU�n��H�V!�a`�)t�W�ws�F?A!`j���!�3�����_7�A�%ѸV�Y�Cdħ��8a�b:*uNu�81A!U��}��J2ꨃߟ�NB7��A�>�`%Q@V���9��g���kF�ڱb0�`떧��}K�|v�JOU���l����:eA�0|y��G&N[�wC�i���ܚ dʨ$�CG4�ɋ^�9o2��I0�s-a�m����}�Ǖ�����Iv����U�GQ��a ��3?g�C�{�9�����z�m-Ԇ�c��;�|2(:߫��P�E��buy���q���I6]�~��˾.Q�7t/xh�x��E��.+`J��MjÅ��4��֟c��`�N1�]�WW\�~\��	�r᪢�44T'$TF�����o��*��`�V��v�W�qd� ��Aķ��ƛ/sI����MX���('V����BCg\/�����N$��f��!�Zu�D)0�`	Q�
Ý	�f�@kV�9D�n��;�KwJ_Oi��W�}�P�5~9�����IPu#)�\��&��"O��_?G��H�'��+!�1/2��Ƶ*7����\���0W)��"��;+�ئ�+ ��+J\W*vT+h����P �=	�߱�֭	���IOyo��A6-=c���ԇƌl�]D�'�}�S$�$�+Rz��
��^{��vdK��Ӛ� e�b]�~�*��Rj02�:�o$'�\Z���}���fbR+"⚃��K��oܷ����2�:_��Z<���1p������"l$4"����؇{��n�����6
c�%�R�'��ֳ���Y��Ɋ5m	�O���9�h��$������9�3�! U�M_ |��m��\'�R5ȏN���^�6����}�U
]%�Њ::\)�<Lc@��Y���z[�4	����܁��6����"t�a��ȲV�%�lV�N���!<"X�y�(����G��Q)�{d�J�q7ߟW¤Qg�X��jF{4}�\��1��Ҧ�+X)"�l#�KK]�On
���5�����aEL�����M�p���;|����P�H��sk ����,3���{>�)f����^$�f$�,"j
hK��?��Zc����������A��3��'�L���Uc�g?|��A�"�?Y �Õn�-g�N�Z؏y�yc~����
����1�T#�`������#k��$�����Q��M�&�����#�d�Hc[��~��!/d��!�%�ec5yjŀ��.I��1�ݰ	J[����J�D��z�a#�Ғ�V~��1,�R���>8)�����0�����֔�/�*�{|h�X���y��ʩ�Ҷ�c �>CZ���5C'�2wN�Hq��7�OcD=�_,1���v�OwT̷qrI�D,�Xg�Oډ<������
W���_�E�P��z.�O�ܥ��������:���( &t�0[kj�������Y��k�(7�͐&J�5Ik�}����!��Z�
�>2�\�(6:y��H����Lzv	����������jq�VuN�SP3�'J�RN^�l�n�hT@b��/��޷��~֜;�@�P�&C�}�w���@`Vv�i;6��!g�����bj�����|&^3��h�-�N	Er�8�B^�B7�eO'��.��~�ç�6wB��&<�R�%Gs�� ?��Z4���i#l�'�g���5KY���
C�&�I���o6{ ���'\2��n�v���fl=�<0����W3��97}��[��2	��� �DNԕ��ٰ`JP]]w�&P��$��sI�b�m��혣az�%�	��	���J�@�j�L�C>���%���9f�o��+q-"m�{�!��_S�%�۴e�O�݅���c5��HϘdtJ�Z���8��n���:~K�� |�6hS74��T������V,��������=��P��R�Z���+v�j�h���F�����s��}�9��|�p	VV�P͝��Rd�RS*�qR9;��2z=%��0Fgt"�' ]�l��#�=&!M�tc���+s� vWL��K�!g8�+�m� �I<I���{U��v�1�hr�y\\�{�|���.��!����?n�=��c���ۚ� .�2����
�]Ӝ�p�| �ˀ+��9��	��LM�����s�����s��Sj�ɓ��{�I򜖸�2 �� �.@'YnG�O�V�'�|��W�k�Ro��6���,�u�5}���ү z�Y���%n�`�y�P����K��+ӬZJ��`�@j���߫ ��|)��z�гJ�����Ƃ��`)L`���%[���]�H���^Q^�n���*h���!�:�E  `ax��������<g����D�t+�&9<v�o���oǬ�*\'4���b�3Vҽ�A;���L����k�+�p������[K�����
��9HO�� �R�"�~�S��	�����F��~�̠�̌N��2~䕃8�:�i�p���Y����JD3����lX�V��S���9+e'��4�i���\��)^t�Y:����̓�x,#�w�+����^�=�Z��0?yk:iKE�Z��חv��ȍ#2�4**�q��M~��p�MY��-��&��}l�mʒկE�`
���9u�����88J�E��_��v����R=[%�!�Z�;�g�rp��(�ؖ�M%���쟥����:e��E"6Ҁ˼�q�z�ق)ɋJ��Ɗ@@�(��P]5�{1�.iED�h
&���*����vQ����Q�%�vB��w��zk
�^v����8��J�5�ێl0�b&����d�m8*�tw��~�.���jzji�ƶ( s���:į���0���f����K��_Bw��L�/�y.�}�6���E_8���S`®�T�����Ne %�#��},��F�.Z?�H�--C�+]�}�t���t�����j��%�e���YB{����k��w��B]���J�4́�%��c��W�s�ˮ��'���9J��҅5L*q�#�}�Y4��n}M�v�SH�������w����X�}f�{Q"����y����U�#�ݦ�|�k�naKEt7W�<�w�������Tm\/�y�ٴ=P���O�<��|�%��4p�vGV%\�oz�`�,��ҿǙ��/U6�a������b�c�<��P�����`bK_5��'��e1/q��GEHP�'"[�E-�Gf� �Z)cP`���c�X{�AX5�ɍ,#S�1%[�/7;�ޒދj�:����≐Y:�"�2h7��t�����t8��k�=6����ox�qa����P�d@�;4i^;���x��{K�*4M%lI�YӫЌuG�0]�:���
6���.�J��)Ǯ�!�V��t��(��{�n[qF��%��8��H�@�"!�ʓB-���s��ǘ/�M3�� s���:|;�&��Sۡ��!��Ɛ�8��*�ĽQސ$��o�$#1��Nf���8�oX(/�+ �<���Iu\����TO+R��2���:�{�¨�8��?M�$3��_�#����_�)�R=%_��pD�Y�YM7��c�FS�e�{=)��O�Ss��=�����#�xB��WOLAn�M+���5K#��~N�9i=v������KD"F�.���k�f�M�G��8�,f��띦�P7�N�M��<W�� }dǚ�m��Ԩ�(R$�Q�`����C����Q�j��BdbRV8����B'�Q�U�ɏ'�Fյ%�7�q5B��e����ֻ�b��fL�"��9�� }g����anਕW��7n�˖t���~�b���F�@(>��\�bX�M�F�``9�m~�h!����f>��� 8�l�|�3����|�yr�N�J���)�v����7��|O[g&��d+-�k�, W�<�����x�U�/��y3�1�re�TU�y��K�:�$�!��I7���4�U�7R�<�ƞ�5�ା1�j��}|���K���4��]BN�$��:�I��n��I���+�cG�xn�f��ي�_B��!|���E��	����T�����8�賡���L�p$u8l�ɼ�U+���1��SW��d��n���*1%c��/�������8�~uG��p(I_��м��|�s�	��=x�,O�m���{%����(Ґ���;�pi��	/�I����|�������ɩ��L0���|���O�/o/u�+��q�����*,�S���ᠨ}�ɚ����D�4�4ਿ2��z�à#�%�5���JJ�Q���W�����F��7���EN��8�Ŋ��P�O�1��}Qi�f�7=c���I���x���F�ހ�>J��/Z�QH3N�@c�L�|�L��,S!��W7��k>��vaՒ�~���ذ�zim�n���M�}��Zv�|�+�Ve7�耸e��S�	�%k��Ew�"K��X�?�M�BB�����mHH�>������=fU�crq��[��$���i��|*}?-h��%RZ�K�
8=&N�F��Ȏ��U��&���1`�,oj$g�sX[VLZ�����1�/憮G�~�`G��U��~��n����xZ�� EL��x��/!4}0T��S�[;-�΅��'!ڣ�O��9�x��K6z��
/[�$L�O������76����5U��_�"o	�aDb��	O*܉��,(7]�n�^fWI�:����,-�uˠ�%�i�Fd]U!���<����zZK	@��]����q�[�*��YYB|����Sa/��\j&���	�+�����<�D��-#J�Bn���4��Y>�[<~�m�*��amx��?���e��TlSc��o��A<�yH�vL�����<�X4��9��$���Vq�(��h�7�i��N��
2�K7f�P˗�?N�G�����-��Eu��9�Y���	O�+֯��B)5�� �5��[q�����mΌ�}|�l#�$�5M���d�9
���Ӌ�u�!��&ۆ݇Mp�E|asF��[XqM��ڡU2z|���ԯ�Z���NS.X`� 5:�$�N�w��`�Fگ���U\�U��s3�pi�7Ƹ��7�\+ #o�J@e/f�Pb2��U[���d���{)���8��.�gbNN�_�{`��\4���F�AGW��-���o�"�r���+��~l(@=������mp��8�zt�:&v�����F�5ּ^Urv�⛪����K>Მ6��ڻ�	M���������X�k�J�g�(�������p������E��uq H��e[�^���2e��J�qϝ�
��1@�*ztخbּ���~�
�do�e�2�X���s}C8Vlе������T�-q*��Х�,��y��e����v�~�$�O�.+�U��>���ԅ9�Ǔ��%$9k+C'�3A����ʴ뫋�j׏��컛+�pN��0�nH�����a�.[)OfA?)|�SL=��R��1�͋�����]���'P�B9�a���ѻ�PO��?�3�	0G���/v́�4�Okщ�AC�"����0�́��9E4���#��\��*��ìi��oN���K嗩����{ŗݜ��d��qe��pG�b��,$�iI�ك-!�<0�׫|�����V��xt������<�,�f��2J/�����������9Ǖp�z��4fU�5"u+��f����ȡ�+V�$M�&����j܎����>�|�oZ�k�6�.5]ޠ�l�m�����aʯ�w0�]~>0e�vEa)��
E5s����֣#_w�)\����CB^,H�&&�OԘ1/>]��홰�(��m�\7M��>qa�H|S+i�I�ivP~vPL�$�\"�i����X�
;4���ԅ��@�q2MVϤ�g�_���(����閂��G D�x:��l������0���� �0����L%��T��D�~#�ڡrNi�X�{��4��˴;X����:{��S�BNf& �`³�Cc�݊yҨ4����I�s},Fdx��5K����R�S�qV�j�VYx��m?�����;h�2Ru-<b�%q��T���&_Ҡ���rӞ���`%7"�h�>�`?�R XR�\ޭ��)��;Р݊������H��H�}&ـ������8�a p��~�$�OSA�{n���v�ކ	�*o���:��]�p�x���:H%wSh�u�~�x������
h}���90�{i�ay��p����!��9���Č�XS�m�g��w�"�� �f�4��1r�W�D	�G�@AbKw�rf���~���Xg4��u'粟�*������b$�����0v��Z�m�b�E��p�};�i�gg��$oO��х�d����ys�y�&�g/�m�C����yl:,�4�ć{�@}�;����.��~\�7�~�!��{=e�`\�ݢ�m:?�fS��3��o�
��E%���GR�}̆;P���^B`
+��'�ɚ��v����{�Y���o�3(Ǒ߸dq��)��L=���l76&̿��Bi���v�����^t��A�g���{���7Xr�,hPM���N���
�B���jƬ}��60��Z����'�gI�,a��N	�-1�qQ��2g�x��3&�h���pp�n�Aw}�%�"�D�.JE-Z���_DH�- u�Ǹ59X�0�q�[]�l��^)`�e�3B�ڎ�$#�ѡݣD��)�4UQg��`�-�'�Q��V�[�E�s��|������vX��q!
�M��(�,�����V�+���'^�'`mQ(6�[l%He`���vd��;Ղ��Y� �`ʋ&sS � �w�ܻH
}F!v���C��Ϣ�6<�)7q�^���o��"2T-�|���W}�ȅ�>U"ZtX+���/�'��m�z6P�/L!	��Q���Q�~�{!TV�6�::�zw�{���[sv?� �`����K�8Ă5`ib�+f#5��cO��o��~Z����H��J.5"娗H7�N�&�����̛m�dz�J9��.WiU�+�ٻ� /e3-=,bv�� :��"w�B^��mP���I�r%*zn{���ٖG0��k�	��![m>�_�����%�S�w?����1�,��j�KP�T�/��P�zN��z�>x�a���p��'�/�Je�{zQ��x����}s�� �/m��w��(N��6 .������6�;��'��|d�����)���!"J.hє�=U�"<W5	~g7c���<ދ|