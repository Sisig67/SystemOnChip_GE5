��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%����!�rr/I���b��ٽ9�K��0�{YYr���o���B���}6��qt!#��-����S�e�QUL�6׀/��,�}C��$�+#G3��U���9��>���N�Q���ۥ׬��8�W�?cFb�?�� ���P��F�2`�7Ll���$��E�eGtA��Kn�:�Ld~�4{9X��y_�l�hNgam���J�N��f��G������kdYr��آ������ϗ񚋻�/wQD� v3�m�)��	kǧr�ό�|*��4��������	Ex���D��r��_I�pNy�(� ߏ��hf^�΂�������Z�����ꡢ�/e���`��,�e�y�7�	��P����	z��5I�"��TG�x�k��%����9���\w�UQ4��-��x�݄LO5
�@B�h̿��b1K���؄�`0��Aճm�g�����8�w���)��y<�m�
���,�K�m_�X�=G*o�&d9ZI��i�-��^�zaZW^l�	M���z�Q���q�e�h�\ԙ�Y�:k~>�m=��[)w�0qwT��$>n�������Y�z�59�ɩ�%�E��r.>�����e�隬U	�����a�S
R��"+o��$�[����Hׅ@.��PP�p�������^��P�\��(%k�����]��WfG��i�ô�1��KӉ�x��^��a �}��[}�dp^҂-:�@9��A�qXkM��?���ޘ����� 5���2�ƣӍ���L7��y��i �V��+?�V�����oo�|g�f�
���z�i�H0X�O�k���@��BYMn�������\`K�Rs��.�8
L���3���G�S��R_�!8vB3�y���o5�?=0�n�B�w}�)��>X���ʰ�}�y`��HZ���'��_��v^��,�[ ?��ˤ=P���%��z��*.���L��C��~���\G�A�y���S�=�͇��Z�KG7S;�@��6�Ro�:I���,�~@;�誻yLEF�7J�K�p~l5d~�븿�Mn#σ�z�z(���s�:xS��8���J;��?O�v��O�a��r�.ot���s�>7��,&�A�%�Li�/��l��S�\P�rRUh�����7RҖ������h�ԣ��O2ҩ�����0�Cs&�!�Fk5W��}b�0لr͚i:�3�m|�ϊ��+�{�&�OeRǦ�鿂�_���lƒ|�f��Br6�)�H��V�ݧ�$
��A��B�V�_�e/�a�"-��3�x��q����CK�d�}lm�77?$�zd�K"�W��֨]#/��/��_����S�KY�j͞���$?z�9���X����S��>��W^��[�bA��X4�1/~v ty8������g���`�������]�0�vܥo�Ժ��ӆ������w�u�(��ԳVh�Z��g�;az���94fN�L����無��;0K�+5&�lӑ��X��8�[�ރ���哽MB��ܯ�D�/�o�F	^�2u�k�]H6Ux�Y�9w(m�������u�Б`j�E"(V�
�o)�c"��o�]�Fب«('D隮�O��,b"�?zɻ}RvJ�WQ�s�~aw�&-�4W����G��d�����O|u7\4��TN���ǅ�+.�ҳ1�^������'O��b���܎�%S�ߒ���1����d����н3�y��^�ak���2�_�q�����'�i��$�>Md����2��ej�6��q�D�l�����C��k!�f^�F�L��0�ӆ�_5Ϥ�.s�)�kſ��ޗ�_@&��2�M��� �>J�v"dD����8�`��/��嵃)��b ��w\`rU]֪�};���J�Kv�jY�F�Z�.p���ڊS�~��Ʃ���2}��u2��&��K��C=�3ٙ,J0�J=)l}�� �7��C�R(���ț\�m[�f-i��6�n�n�(�Zw3��V_�N���j�|_�g����pE��j�׌��Y��ܛ�w	�j�D=�h�	s�C�L�U�x�e��0���|ҷ�N`�x��v����U��oFڀ0�K��i��m-�<��jZP��zT�	�x����AeFp��:<)JM�-���~�xlf0���۪tydA��C�A��N��oL��9��fT�w��Oh
��B���r=�q(�kqc[�;(#�jW�&DW1���	�XOԻ��+a��z�&�^b��f	hq��K���~ݰ �gƘ,Z��`Z.� ��҈ޕd����i[�V���m��2V�?�Wx����&S�����je��Ip�r/�'��.tQ����Z�\�|���%i������H;|3�'�z��)��S������8���ΌE��xp1��Vũv����ĩ�k������ҹ����'m[}n�o���A��!�w�x�@�xO&�	�=9Y�q͜!���P��[tiٻ
��Y���
��u��V�z����.Ob�F68�-�<�KI*Z�$�~�$�*:�ăG�ब�:e� &�Q�<�S�ݟ
v8��*�1�?�_����k?JA����U�m�}�K(���=���l%����5T�
��SdS���$��o,	u���s�ծi�h���|�(i��T�:c�(�!5�f��:.k��H��5֎��O3�TgI'O��QN��-�א��+ӗ�<��UEX�ˎ9���}!�F��K��%�I��>�8���I({~�6���vn�V9*T�8ȉ`z�06�2���r�m��$��~y��$	U�fhp���l!����Z&�!u�]��n��v*�H_�[ �b��oj���<�<0?]�K��`�ǽ)��������̀nqS�h*Q�h��X�y*�Qk�,%g��/F�6�q=L��;4��I��+h"�@Y�ֶڗ���~��c\��N�",�ψ]��������a I�S*��c|BS�^�������o{�]��w��J]njr�z���0=G��I<�:<1�M*�-����&¢3���KG7\K:٫/�cnq\ZB8K�|W��&3ѝ ���en�]�;z[�%�{�_Y#<mꭞ���� 5I�S�#�\.:Ѣ���}Tu�Gn* �6��P�`��Ӣ�c�A���.,9c���וֹ��������m��E@F��$jK[���αt��VaPk~B?�t�a�ql�*�$�8\W��J�.���D�I�FY A�I��F��/P]= ّ)Ű�;RT�%�o���@j
D��p�y��_"8N+�P��	�<]��r��nUѪ8C����ǌ�ʹ�6�,���� 4�
��m���N,=xR��K�\">�E*�AFj�ZĐ|s?~�'`�O��N�U3^u(����9�+/�}bŮ�!s<���^q������.c��0�xR�C�"�Au�-�b\o,l��V��Z��~0�c��E��;*���`N)i�w6���'��\���g�l�'>�B�cB3����5�ICDҕ��z雫X����X��w��!���;��2^���U4�Z}� ~��3?�쉇�e�.�1�.£A�O����g��� �"H��u��"����C[�C} �㼔e�rjeP�S�V�������M��T��ώJ��K�(��X.��,?�cӨ)��FY����p�s��y��IX����em�����M�B�W[��)b��N>�vi���M�d��W$V���=�a YR�N}�W��h�>.�Af�kq�Ԣ��mK;����2���S�U{��Hwg�gD�1�īE�R��Fjl.A���O�jq�%�3��v����o*m���>��0Ђ$��i)�V�̗�wܥg���I�M�8-�������	��񜞳9���W�J��`�#Jk�R�{�g`
�
5���f/�z�8�CSm°2H7R�<���������G��-|~E�q�=����ȃ\L�sN5�E��E���5�M��T��M�ߵ+�Ik	�@��ۺ���d-�o�ar��-E� w�v��\�\��y�DA�@��&_�S��/���xIm�����}��U'$Cc&���B�r�����U���~��z��/�ǉ�_�<i*!��Ŗt�����c��Ϊ�p?�>nQR��Kc�5�������ɞ ��Q�Az�}}9ɒBЌԷA����jrCb�N�Ae,s>��v���`R�J����Y�Xp�O�m<��53?�|R:��xИ�R�E�C�6��h����T��:�eƨ�Da�� �:O��5���`�og�T"C4ތ/F5%E�������\��ʽC��#�(d���)"κ�W��W_?Waz­�fr�*|P��:��c9�9��ۥlO�9�� �g��J���a߰Y����̼��N�u.Bˁ����T�hm"#�D'^4g��Б[h��~-�ߠ�M�������դ�0��A2��?u��Z�Qm�+�j�� n����
(*sC�2��N�6���2�v�9홓|�Gn�	L.��&��s�{|F�qRrl�qV�=x>/���_�����c�A�{`�t�ق"SA(V���l���RKT���~g��L�阘f����]������Em����E��B�tZF/n-*�ܖ������OJteʾğq`'3�p�5��9��^�y�ܢ��;��㕄[k���6�����ܤ6��WTe��gq*�o��|o�vn��	�Tg�00]��o<n�	�l��R�� �W�٦�"[�>[m;k����]�'��Eʦ�&�8��G���T�b
�L�.�o�L�z.@�4�wy1����(I*`6йHE��F�->�`=�*HP�I[�	�l<�sl�<�O,��v
���R��߆O�u�p�����rB�Q�����&,�1�,��?r�]n5�i���+0p�ҵ\�w�nG/��^C���\��Wީ��6c�8f��Ӧ��A�_�		����Πl�q����1�h�'��璧�x���.)�Z������o�.��'��BHS��p����{O��,�����S������	�9�Ґ�т�/�p���[��u�U���
e���8�G֗J��Q�wP<�7Ǡ߮\F���D�Z���q&����E{�gOX�V��CEU�"/ux��Ţ<������u�ї��TB�\�=����#ŝs����ke���p]�v�%���4�:���Yɽ�w�5��۰��=��F�'�m��/�ȀFu?�ҫ_�7VO�B��mo-3�E3D)U)ļf�5�}0%Dr�+y\>\~i��]U6�ڻ8��'�T��_�����X�I6��B�LK�4�>31p#�'��A{��q+�u�����a��:D	|�66Qؑ
�'3��.q;�7��-�|	��ͭ�\X���隤J�]�������$y8�|��;BJ��E�>�q:���A��)�FQ��s���}�:���
��@>���:���@��R;�q (�e3o��p�]de��i�X(��z�C��eo�m�u�e��#K�����*͟b�.����*�ћ�H�q�b�M#�"�y(d��}'�Օ�p�r=g��>]�)��_�~��@�#�p	�U�h�e�g��!<��G��kL5_]=����
��j�|w�H7�3�7*���g�⡪��
����PV0���W>�������R�X]<�;r�P����K�-$ƕs����x�J�c�ϥ �U*�4��:�BJ���8�Q�7�a�E��54�Ͷt[�%��3�Ԣ��*B֨��5lr�t�(a�ϊ>\!�SA��/�Ά���/z��r
��)X�|3d �I��9<f3>�'���i�f�U�%CI F�aQkd$Y��'S� ȲXp�:#�풏��|C���X*9�Jt|�&��| ���T�s�Mѧ�l��"%�i�e�7�2�����R��]�~���7a�A�xA��焮v�-T
+�f���?�ƟM9��c�ݓ�$�U��F���F����ў:�G�_�P�P�.�8�h�vg-�{-/��&[���?x"�J���8W��J"j>9?I�2��-utn�`Ȟ���%��܉ku4�?��37���Z���ln�E�������D�wɨ���zZ��R��J����۴��^��|!�op2����J�+����Aq�%�%�z-�%W�MhX��=�����y�}���M��t�%a]�N*\/Mb]W!��N>}r��{�.�bӱ(�c�)T�ң �zIP�R��T_R���)�uDM�#YSŦ����J�X��خvb:3��hw2?�3���+��F{O����c�I$E�P`l��T1���.���K�!�*��|!��(P�X���9���ٟ8^e��C��-n�=|���o�rⓡ����|L��$�%�v��wYD�PЋ�����F�25\E~�k��{#�I{�d��o�3����9-~�*�=&�wK��;\ w~M����󇪁��<���ꔿD�����>��Z��Q�Y(�9C�g׆n���RV�5�y�#��~���"m�@�� j�^6�d��u��1��A��_[%LpKȨg��>RL���-⤟Y>p�k#��~�T�6og������'��LZa�S/lM�V�IZ��ʥ��m�r����~���; 4٩���=��en;��+�$+8��<D�_�7`)��7ʩ�����j^���R���;4Ci��ZЀA-�O`����������l��|@M_?���I�'�uy����o�e�[�[��
5q�I+�D�	ޗ#�o