��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%��)��/H��s�<�8-	��,x��9z#�T#��`�A���n�<��#"VJ������fWs�5��+�[��~#�ۣ&�u�e����J �@��O�3e��ėݎ�i�yu�4��nWU�C�X�^��HC�����_<�PPb�s)I���W����=ª.>�1��3##���T���oQF�O/����­32eD�a,s(��A�*���K�����$g���`��d.G	�D����
)2�����J�;��
�௟B���-St�1�n,ۣK|F�b.4�����!�nƦ��p=��˔}ϭy��W��3Hꋃ�F7��QV�o�".L:_�T�*�4�U�}�FS�jR�U�Nf�$MDF2�L���U	�؞"�.��&�I$�Բ�0G�"P����bե&U��t��g���G�DJ%pN���9s���Ãx�3��+��H�١z���oH۸��\t;��c�>��I�d$���iH^�'��E{˰�|�$`�\8��?�Cc�P����n�-�J��>�a�}�k}H�O�{�F�����!�0��(��إu�A��,�[��	_�����^��u[N˟��� �92^\����[E�P�u�g���x���]>���oZ��@�#�)�bMI1o]ٖ�x��̆o�x8g�=/�ם���0Z�2;���\�a�mU���|���e�¥L��BSsbߊL����RS�3T�����/���Z���!~ c}�-��W�j��|~T��V�7OZL8v�f����J?J ZiU�_��s�N6h��yF$x���7��s��=�ؑh_86�w�����R�������mu���P7ຫ^ a,Me��!"���ډаx�)?Ŀ��ˢ��j��1@�wU�Kӎ	~p}�O�J���#X�ѳo�2�C2>S�ŵw���z���)H�Z�z��U1z���G�~�O���a�'��?pliP˖D��M?��!�� ;������>�;)
����������C=�+W�0���w][K�0��G ���-��2qj����{��^Дm�
KjT}�1�)�5��_\��*uM5�?� w�����)��/�ST�b#�/�:[��'e_���R�Z�`������FF-�?U�Q�!����8RT�r/k?ݨ��[��M���2/l0x����ǖ�ڢ�;W����A?*t�Q0塏(ۏ@�]C��^���Р�����:�b�v�}H�qb
ם_=�R�H���d��3���6�*i�(�gWb��hV8
1kA
���uE��1���)8[�;t=6�p��j�9����'�Ry��L2z��:�g	 �"{���.z��|�z���\[�m31��@v�N�c�c<�!c�=��%�o�o���'�? �}a'�"pĨ�A�����Av{_F�<(
��3y�ȏF���!���*���n�;w2΄�L�X�L}c2R�IN��e�QZä��sݼ^vI��|����G�:�%������#�r����n��x~���@��ڹ����/��&��!�'�Y�M���HHM	U=*�T��cu���O�곿 ���쌂��W�vOb�}�ٶ��TH tא;|��@��x��KSHچ��FP�^!����:�*m�N���`�>��(Jl��7x[�b���(��A���ѭp�8�c�p�IU���^�D|
=�f5=��5�T4ErR��[�'ď�{��']��g=p��J���S���jwF����U;s���~�#�5Sx��#��ɨ��@���t��^*.|jb`P�7�r%���E����s�z�C��Pߧ/gd� ]�쯯�S���1��d�5S�
��j^�6��&���'q�A�s�@���aq|������Vj���;�f[k��#����qo]�*�'J�� gf���U�o�����#�^X���#��G��yp�,G�={y<�3���NC��0���ȑ������ �w>��(_T�놥��u�z]�7̈́�=�M���#����[]�ֹ��b���[P�`����+�9�ߒ�+.fa�ͥȞs	�H���|-�M70�����މ{xL�/	6$�MRN`��$Y1�  ��/�l�Z:���|��S�#hU�h������{A��O^��"�1f�ʐ��G��BQ��,|�D���?�5h���Բ��̎wU�9��4�'�ty&�j/�Z��������5�J#ɝ5�G$m+x"�`d��j������}񤝕����f�)!J��O������s�c���"2���5k׍d`��:����݉���!5H5�8�,C)�f�uͬz����!�� ���vcLCslް2ӻ��bO^�8C|r"��S ���q�ԷUvK�	]'�����	�B�|�\���We ��IУ�AG|���v@����h��P3��B`.QW��AcS�S��S�[�� XLI-��t� i�S-�x:����e6�t|ȁ�ۉY��<��`�C@knB
��zϠV���$P<;���ek��64�H����AYk��p�,�ZCZ��B�x�|J�\���Qٹ(�o�Z���8����W_�f�:�d����a�R�@���p2��Ea�dfY�bm�H�(���aRP����SI؞�%��.��Mm�ȏrȍ���M�N�m�T�}��R�2[�s��F'8�tOv(ϻع �����Sh��_�ǟ	�� ��yW�r<�Ȇ�A!��m�%#\�*�
[#��gt�
`h ��;�j��@�=f�(]�:���as���^�|�Ӑ��c�p���P�K���/�.����J�,�/8�^�F0��l�!F[�ۢu�Zx�Qv�;�f��dy@���R�տ߫�xo\�DZpX�|�L�c���ո�"7��cː�G�Dd�U�q��
�_'�� �ȟ����b۳�<~$4_�h����?��h')�z7�� HhDF����?q�pyw�8�̒��ll��}#o���)f�|�0�` M5�&R-�{�z�Bե��l|5}븟u��,�)C���)��&�N�˫�0[=Q���_�:��+R�򻭴��y���	H%�G���fZO�L�c�%�F��F"�0s�~NN�����R[�9[���E
kCR3d~�l
s�Ds���:1u��Š���?�&��<�b�ÈzS{k�;ه�:U�r����RI�y���	+���Q�&2L2�S��D4���'۷�m�\Ǩ�
"#]m�[��A&z�"���!���5C�����|���r^Vg��>K�6� W�h��$����R]k��T�:��=*٨[�<�����i�`#�c�P����iΈ��ں���h/�P��� ף�e��^ZO�*7hSױ�\}���>z����,k8"M?`��iD&�<_�@�� y��ow$d�TT���)T��sc���e�|P�ݳ�&M*緶�ڙ��b���ת��֚��g�����ф��ӽ[r�U��K1��@2�G|B�-�W�|Qh��\w��=����h�^�6S�W����D�I�� �4��Fpr��{8���v�_]e5���(��+�&�mv1^�V�䶔P��Pm���}����e;������M������ϱ�z ��^Ԕ��"��mq� Zԝ�}���|�~�-�sa*�k�l,�C�6}���]eY�z�q�W��arN#f��J��Z�<��7�`�u+�Mr�E����lXʁ��"yE����Qu%��*͹k?�Z�����U�qK���κp��Y�D�T�WEK�*JX���\b�v�|��	ܲ
�%�}]�B��/�J�dΉ,2���=�R��[=!ۤ�%��%Q�oVL�~��=�N̑h�UGO��R�Z��K�����%��<ty��Xu=xW4�`�-��qխ�E�py�C .�c.��A;\�ѠTx&	�pw�{��!��� {q&�l��������5'�"րt��.qu+�C���X8�;��x��J��Y��q��m������۶	MH�d$�}�ȸHp�6�F���DW���w5�}�P����zmXo�	S�P�l/^i_h�0\]���??�	'�Ǒc��w�i�4Ub�
����ǈ�J"�[�8�R���}o��g���1��|���-�g�.���Q��u"�W���u4��!�Ӄw�p��27���Կ���Yg�	���7-~���@�?r�pG9eS���@�� x�^FҴ
E��P��2�n���3����JW`��T�Ίx��rK�U�Z�c#,�kNi�����h��T�q��D�dv���$� �ޝ���DA&�7���a������)s{N��w[ O���䔭�
��qiV�/u�E���+������G�+`_`�* WKҧ*���?��2,�)�2<�7��d¼��-�9(h}%+�_��X�