��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj�o�v{'����!���J�qL�h�5�$a�����߀���9Է��a�1 g9^r�M��*��.ө[?G�G(�wYg2FZ���*�Ǟ+�	[rt���C��E�z��r�X����cp\X��;�W��
�,TMW�6ɩ�p��&�1H0�o�'��
���.tP����};�y�.5Ȱ�3 �Ղ����y��G�A�?��\]��h��V{w�ny~��p7M(�g�Jߌ�a���6K�b'n	1�4�5���؈��IE���,|���Ac�1O3HH�d�8)��1"JY���7	�QI8����I&)`3������#��-��p<�g�)Q�g��ė@�:y�'�ٱ>�~��y���!�P-M��̲#k<�Ĵ��'��r�7T(�|�����Ɓ��&#�P۱�P�) Q�8WG�ˏ�@ʺ��H|��L����̑������Tx�!�z�3�m9Ѣ�{��5x�^��Ҹ�ځ��)�[3O��^i�~�����ߦ����ى}ڛ�a��f|ЌaL4{�r"V��Ġ�g�bጔ�t7ۮ4�nlr�׷�rr�F^�9�p^8La�Q0T�,���Eak��� ��V2�Ѕĥ�fqȖ�1},���� ����V=�'A��@�x0��|�>�zdT��N��0����4��-9׹�g����&�gN^��{*�&F�N�l�{�o&�ۘP�����N�$��Ā��~����$����^vH,�nߞ�zCS�N�X�u0�x\W�c39�ϖL�3����nOy^oI�.������vj1;�9�F��j�!�RU[���B��Ap�^�>�$� cZ����ɜ���
�,�ܳ:�h�j��Oĵ�Ik���
;`���%�>�I�E����S�IݰN�`jL�·��cJ�G-�:�z��,�NҶ��@H݊������W�