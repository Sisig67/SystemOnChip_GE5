��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%��Xh|Rk���0�Fg�������3;E�:��*$��΂m�;�2L��ݣ���s.x�`���@ý6�$8xQ ��m\�1������=#1���*:k��H�H�Z&�s6��-`�3��ʅf���us�Ľ��S�U��yEF�t���� Ag��1�*k�W�X��P���R�~o�������4�����b�*�Rz���Mn/��b_��k�w��wu\��z���cS�t!��%
@p���V�h�����cy�	i����^ocD��ڹ������ $%�k�Nmv'OOH�Jݏ:�)MI�X��Ճ�J��۵��b����@�mM��e���_�[��76��?U.�W:�/�S������<+��"��rI��\q��,�3�a{]�º�z�q=��g!��@;��R�����i��e.%\}�PY�V1��0g҅(W�3#{��N�Mn�*C�j��?`XUti4��˄�G�w#.
� ט��!!�O�	c�2��6P�3H�,��LH���j�=�����A	{��F�AA�Rm�� ��$`D��n��h��E����K���&�����$��~���ڰ0���PK�	`Ӈg_�a��9���+�7����G5!���~{On�!坝&�?_�
���(��Y멯�S�A�9�� �w_��9"�z7 /����≍����x��<�&�:�tK��L<y�}����ȃ��f3�NGyz	>���g�X�vՕ��������S�!�w���z ((v���,�߽X�cb�C�yLS` �P]y�vY�,�������1?�fH	V�F{у����RR7?R��o�H��8�� ���0RV-e�P��6~1�9�SyIʿoL�ʹ�G��Bo�4
��Ic������N2N�i_�j/$/�(u���$��2nY,��&q�P f������DQL�[q�$O6VN��7�v}�襵Hm��f�x��nsnΘXnxW^�I���<`{e�+M��t&�KU�d�ƿ�UΈ���F�B[u����ю����ӳa0�`��[a����H��d�ۛCf�}p�����.��5hs�������l�Z� ������g�J���2:VǷ�V�ƒ���j�:�fG0�@�k��#Av|T���#$MHc�i�q���_(rI����'hTk�n�6��~[���JWuC.0?��7���o���g'Eo$Ʒ�F|eF�1P%i���9�y���g��y���y�|�EA;����QX�0��X�y�/8��VW�(��͢$���]e�>�m���[;`�����؆�Kw��D[�-|�U~���M9/><Y��~D?�{*<�(�5~�w�z�f����&�����J"��~��)�0k,�@�� �� +��}<oy���Q��X��P�=Ŵ���ew��_�RU��V�WH�"��[+Z�[�~�3J<*�^����&���P<��p��~���s�����O�k�Dr,&F��� i�=�2P:��]�Q�U;|D͌�^5}��w8�":Ð��2�&a�cu�`\!�����u�Zӯ=�R�>i����SF�@1"�y�����78$ndi�����]H1D<�J�H7"lb�S]b`���r���(K_6���qC�|�P�4���jη��������Է9����(p+��]�ƥ�yQp\�M�',|O��b����f^��"��2����DA5xM��H	��'{�� }Y�v��R2���d�.09q�F�q���b�{��L%��uXQ����x�5�%G	�w�q,bk9�&�x���/�h�������+Ċ����;�\��3
��d����R�z7!��4�6��)}:�nJ�Z� �E �����oef@0�a�8��C�s���9�z��q�ЮM�1�l�~d�k��	�ͺ:��m�e�ձ����7��N��m��k���g���	9P-���&łh��qI�^��	��"���8�h�*��sG�n0(Gt��s��� ��Q��&0�Դ����utN�Mb�ߜx���j�G.��F~��1#�.c�gG��4�"��0)1y��SNt`\���ZM�0$��s���V:�Z$�Ʌ����Y�&���[�v��Ģ�%>�-����;�����!�q|��,xG���D��xvv��wj�3)X�����a Q���1�q�w�]�>|5��02���6�T@���!���_�Զ�
`��2s[���dJ�=���|�˓�Wq��d���>��X|�v
LC�o�m�ᭌɀ%��������h���ֲ�>N)���_���y�6���2���ۈ���B42�5�u�KC�[��h���ȃA`R*�k_����]�V����`��Y��B�@�ei]��k��ƨI�u{k1\�2ڽ�:�}`����Nj��7|���0]��O:���z���+%�4�	��������C�3����[h�P|��%� �Wغz�wX��2��Yͳ��),�������O\�V#�E���z��4}���%�;/W>݋���&�iF���Ju����'E�;,aʩ��'��ML	 A�>��C�Po�?��Q�?^hެ��]��O�sDl�gh�짊U�Y9'k���7T��8���"%��Z��ܴrcTU��T��QM�����*v^��
���N���nZ��M�G�	��q���-7��X^�\�ä*L;�hc'���R	<Ŷ�_���W41X����X+���k$g3��(	�-e������+C��l�����%🲯��B�~������w�B��r$ܝj���b���J~����7{W-ȉ���/�I�3RSƦ$"zY�	���YkZFԱЬٚ�pz4�z�@�k��;�tݦ�Y��[6���5Ƈ��&�W]6�,c �I=�&R��ی��UńQ/U�z{�0�?Dk;�4�[�q��m�+
o�p2y�G'�6��o���A�t&��`�W�O7�O��0lb�*�,-'&��<�)�����n�Aj�µ-`b�o�A�.h;)b8���u�u-�w��f�{��ooq�ˬ��W��"Eǳ��VK�j����z���r�/T�Z��W��/�a3s2�u$�Bo>�cbG�uг�8LG��¼�ۜ~%��Gӱ:�����^--��vS�7��s��{Fq�,�
m��U	0w����8�y���H�W,��5+�\��<�Vj�{� �$*�I9'�4<\�6�o�������ߵ������rTjh��R) ��TM�Q�u܋(�KsKU�������"t����a�C��\�b��t�q��x9�C_�w��T;���*j����P�D�9;��&�0,Ob3��)aKG �vgQ�W�}lWrż>h`�(�8o`�`-'~�k2k��$!�8��.�?���:ӷ3�'�<��y��s���y>��y�m�uL��V,X���L�#��a�v�t�#�Og;&�<��P���Du�f�A k���!���X���ژ?"���ܟ~�`�iyPv�G߁�*2�li$}8�J���I�?"7�iQ��ث7��e�\r�n*,�U������5�{�>���l4��E�蝌M��W�� ��g'�7�?��\퀠v��o��eX�Ҡ#��3�K �	��1z���d}�6�N��Dy4�����h�͸����RE��K��3l�z�C�8^������"�u�j(�D �rޢ���Tڙ�=�"�Tq��S[�2+e_�DA�u����c7� ����
?l�>��v�X8�?�@o{�����72�RY�9�w�����K@�к����xګX��c�M�"�k&,�<v<�4���1���@�%��\�@�ڦS9�"JU6��ȣT�r�J4k�Z �/yxՏUU#c�7�=��L�8������,"�M� �%�KLѽ����ҟt�
ؒT4��=���{�8���ߟ/�6��s�{��eʘ�=�'\�ʂ+ׄ0d��ޑ��L�?c��S�
��b��]p��{?Z�`����*�XNZ�7H�u[6R��yFg�p�����z�֧C��K!�����x+I��)�p"MKi"\�[V�]�x.x� ��f�|X���) �%���3��R�L�V�	.�`)6$ [2���Њ�Y�"�֭�� ��Ohp�"�� ��L�H�rE,À�l��\5cxoO6�ΈH�𮋇�r�Nͨ~!�������;b7����p�a�2�������5�-�|�z��+W�63�T�[�����S'ٶ[�@jz��L�>���۵���)���?�N��?T�5+������w�X�̮gjS�J\!�ў�6�r���h��^���t"���!�=����tc�c���]:ʥ����Rz��)�n�q�����![����rNp��l.�q�1�����!
^����M��C�cpF�|DB~��S���0��%��54	�����=Ze@���;&�B���)���v+�LT�j�D��}�1���t�2z���V+�4�t�Iz���؉ށᇀ��誄� ����7F������a��7I�B��]v$Z��B�۪mUK�Uc����2MlL}���8�Kt��o��Ca�BHa�}��궸[�Ց`ӌ�O���+է�cƵ2~���u��LN��x��W��hs��W�vt>�����	�rŗ��B�w�`�.�Q241[&G(����[?˔P�9