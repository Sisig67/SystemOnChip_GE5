-- NIOS_RFS2.vhd

-- Generated using ACDS version 24.1 1077

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NIOS_RFS2 is
	port (
		bt0_export                        : in    std_logic                     := '0';             --                       bt0.export
		clk_100_in_clk_clk                : in    std_logic                     := '0';             --            clk_100_in_clk.clk
		clk_50_in_clk_clk                 : in    std_logic                     := '0';             --             clk_50_in_clk.clk
		i2c_scl_pad_io                    : inout std_logic                     := '0';             --                       i2c.scl_pad_io
		i2c_sda_pad_io                    : inout std_logic                     := '0';             --                          .sda_pad_io
		led_nios_export                   : out   std_logic_vector(9 downto 0);                     --                  led_nios.export
		reset_bridge_100_in_reset_reset_n : in    std_logic                     := '0';             -- reset_bridge_100_in_reset.reset_n
		reset_bridge_50_in_reset_reset_n  : in    std_logic                     := '0';             --  reset_bridge_50_in_reset.reset_n
		rh_temp_drdy_export               : in    std_logic                     := '0';             --              rh_temp_drdy.export
		sdram_addr                        : out   std_logic_vector(12 downto 0);                    --                     sdram.addr
		sdram_ba                          : out   std_logic_vector(1 downto 0);                     --                          .ba
		sdram_cas_n                       : out   std_logic;                                        --                          .cas_n
		sdram_cke                         : out   std_logic;                                        --                          .cke
		sdram_cs_n                        : out   std_logic;                                        --                          .cs_n
		sdram_dq                          : inout std_logic_vector(15 downto 0) := (others => '0'); --                          .dq
		sdram_dqm                         : out   std_logic_vector(1 downto 0);                     --                          .dqm
		sdram_ras_n                       : out   std_logic;                                        --                          .ras_n
		sdram_we_n                        : out   std_logic                                         --                          .we_n
	);
end entity NIOS_RFS2;

architecture rtl of NIOS_RFS2 is
	component NIOS_RFS2_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component NIOS_RFS2_SDRAM;

	component NIOS_RFS2_bt0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOS_RFS2_bt0;

	component i2c_opencores is
		port (
			wb_clk_i   : in    std_logic                    := 'X';             -- clk
			wb_rst_i   : in    std_logic                    := 'X';             -- reset
			scl_pad_io : inout std_logic                    := 'X';             -- export
			sda_pad_io : inout std_logic                    := 'X';             -- export
			wb_adr_i   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			wb_dat_i   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o   : out   std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i    : in    std_logic                    := 'X';             -- write
			wb_stb_i   : in    std_logic                    := 'X';             -- chipselect
			wb_ack_o   : out   std_logic;                                       -- waitrequest_n
			wb_inta_o  : out   std_logic                                        -- irq
		);
	end component i2c_opencores;

	component NIOS_RFS2_intel_niosv_g_0 is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset_reset                  : in  std_logic                     := 'X';             -- reset
			instruction_manager_awsize   : out std_logic_vector(2 downto 0);                     -- awsize
			instruction_manager_awlen    : out std_logic_vector(7 downto 0);                     -- awlen
			instruction_manager_awburst  : out std_logic_vector(1 downto 0);                     -- awburst
			instruction_manager_wlast    : out std_logic;                                        -- wlast
			instruction_manager_arsize   : out std_logic_vector(2 downto 0);                     -- arsize
			instruction_manager_arlen    : out std_logic_vector(7 downto 0);                     -- arlen
			instruction_manager_arburst  : out std_logic_vector(1 downto 0);                     -- arburst
			instruction_manager_rlast    : in  std_logic                     := 'X';             -- rlast
			instruction_manager_awaddr   : out std_logic_vector(31 downto 0);                    -- awaddr
			instruction_manager_awprot   : out std_logic_vector(2 downto 0);                     -- awprot
			instruction_manager_awvalid  : out std_logic;                                        -- awvalid
			instruction_manager_awready  : in  std_logic                     := 'X';             -- awready
			instruction_manager_wdata    : out std_logic_vector(31 downto 0);                    -- wdata
			instruction_manager_wstrb    : out std_logic_vector(3 downto 0);                     -- wstrb
			instruction_manager_wvalid   : out std_logic;                                        -- wvalid
			instruction_manager_wready   : in  std_logic                     := 'X';             -- wready
			instruction_manager_bresp    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			instruction_manager_bvalid   : in  std_logic                     := 'X';             -- bvalid
			instruction_manager_bready   : out std_logic;                                        -- bready
			instruction_manager_araddr   : out std_logic_vector(31 downto 0);                    -- araddr
			instruction_manager_arprot   : out std_logic_vector(2 downto 0);                     -- arprot
			instruction_manager_arvalid  : out std_logic;                                        -- arvalid
			instruction_manager_arready  : in  std_logic                     := 'X';             -- arready
			instruction_manager_rdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			instruction_manager_rresp    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			instruction_manager_rvalid   : in  std_logic                     := 'X';             -- rvalid
			instruction_manager_rready   : out std_logic;                                        -- rready
			data_manager_awsize          : out std_logic_vector(2 downto 0);                     -- awsize
			data_manager_awlen           : out std_logic_vector(7 downto 0);                     -- awlen
			data_manager_wlast           : out std_logic;                                        -- wlast
			data_manager_arsize          : out std_logic_vector(2 downto 0);                     -- arsize
			data_manager_arlen           : out std_logic_vector(7 downto 0);                     -- arlen
			data_manager_rlast           : in  std_logic                     := 'X';             -- rlast
			data_manager_awaddr          : out std_logic_vector(31 downto 0);                    -- awaddr
			data_manager_awprot          : out std_logic_vector(2 downto 0);                     -- awprot
			data_manager_awvalid         : out std_logic;                                        -- awvalid
			data_manager_awready         : in  std_logic                     := 'X';             -- awready
			data_manager_wdata           : out std_logic_vector(31 downto 0);                    -- wdata
			data_manager_wstrb           : out std_logic_vector(3 downto 0);                     -- wstrb
			data_manager_wvalid          : out std_logic;                                        -- wvalid
			data_manager_wready          : in  std_logic                     := 'X';             -- wready
			data_manager_bresp           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			data_manager_bvalid          : in  std_logic                     := 'X';             -- bvalid
			data_manager_bready          : out std_logic;                                        -- bready
			data_manager_araddr          : out std_logic_vector(31 downto 0);                    -- araddr
			data_manager_arprot          : out std_logic_vector(2 downto 0);                     -- arprot
			data_manager_arvalid         : out std_logic;                                        -- arvalid
			data_manager_arready         : in  std_logic                     := 'X';             -- arready
			data_manager_rdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			data_manager_rresp           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			data_manager_rvalid          : in  std_logic                     := 'X';             -- rvalid
			data_manager_rready          : out std_logic;                                        -- rready
			platform_irq_rx_irq          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- irq
			ndm_reset_in_reset           : in  std_logic                     := 'X';             -- reset
			timer_sw_agent_address       : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			timer_sw_agent_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			timer_sw_agent_read          : in  std_logic                     := 'X';             -- read
			timer_sw_agent_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			timer_sw_agent_write         : in  std_logic                     := 'X';             -- write
			timer_sw_agent_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			timer_sw_agent_waitrequest   : out std_logic;                                        -- waitrequest
			timer_sw_agent_readdatavalid : out std_logic;                                        -- readdatavalid
			dm_agent_address             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			dm_agent_read                : in  std_logic                     := 'X';             -- read
			dm_agent_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			dm_agent_write               : in  std_logic                     := 'X';             -- write
			dm_agent_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dm_agent_waitrequest         : out std_logic;                                        -- waitrequest
			dm_agent_readdatavalid       : out std_logic;                                        -- readdatavalid
			dbg_reset_out_reset          : out std_logic                                         -- reset
		);
	end component NIOS_RFS2_intel_niosv_g_0;

	component altera_avalon_jtag_uart is
		generic (
			readBufferDepth            : integer := 64;
			readIRQThreshold           : integer := 8;
			useRegistersForReadBuffer  : boolean := false;
			useRegistersForWriteBuffer : boolean := false;
			writeBufferDepth           : integer := 64;
			writeIRQThreshold          : integer := 8;
			printingMethod             : boolean := false;
			FIFO_WIDTH                 : integer := 8;
			WR_WIDTHU                  : integer := 0;
			RD_WIDTHU                  : integer := 0;
			write_le                   : string  := """ON""";
			read_le                    : string  := """ON""";
			HEX_WRITE_DEPTH_STR        : integer := 64;
			HEX_READ_DEPTH_STR         : integer := 64;
			legacySignalAllow          : boolean := true
		);
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component altera_avalon_jtag_uart;

	component NIOS_RFS2_led0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component NIOS_RFS2_led0;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(25 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(25 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component NIOS_RFS2_ram_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component NIOS_RFS2_ram_0;

	component NIOS_RFS2_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component NIOS_RFS2_sysid_qsys_0;

	component NIOS_RFS2_mm_interconnect_0 is
		port (
			intel_niosv_g_0_data_manager_awaddr               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			intel_niosv_g_0_data_manager_awlen                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- awlen
			intel_niosv_g_0_data_manager_awsize               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			intel_niosv_g_0_data_manager_awprot               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			intel_niosv_g_0_data_manager_awvalid              : in  std_logic                     := 'X';             -- awvalid
			intel_niosv_g_0_data_manager_awready              : out std_logic;                                        -- awready
			intel_niosv_g_0_data_manager_wdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			intel_niosv_g_0_data_manager_wstrb                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			intel_niosv_g_0_data_manager_wlast                : in  std_logic                     := 'X';             -- wlast
			intel_niosv_g_0_data_manager_wvalid               : in  std_logic                     := 'X';             -- wvalid
			intel_niosv_g_0_data_manager_wready               : out std_logic;                                        -- wready
			intel_niosv_g_0_data_manager_bresp                : out std_logic_vector(1 downto 0);                     -- bresp
			intel_niosv_g_0_data_manager_bvalid               : out std_logic;                                        -- bvalid
			intel_niosv_g_0_data_manager_bready               : in  std_logic                     := 'X';             -- bready
			intel_niosv_g_0_data_manager_araddr               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			intel_niosv_g_0_data_manager_arlen                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- arlen
			intel_niosv_g_0_data_manager_arsize               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			intel_niosv_g_0_data_manager_arprot               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			intel_niosv_g_0_data_manager_arvalid              : in  std_logic                     := 'X';             -- arvalid
			intel_niosv_g_0_data_manager_arready              : out std_logic;                                        -- arready
			intel_niosv_g_0_data_manager_rdata                : out std_logic_vector(31 downto 0);                    -- rdata
			intel_niosv_g_0_data_manager_rresp                : out std_logic_vector(1 downto 0);                     -- rresp
			intel_niosv_g_0_data_manager_rlast                : out std_logic;                                        -- rlast
			intel_niosv_g_0_data_manager_rvalid               : out std_logic;                                        -- rvalid
			intel_niosv_g_0_data_manager_rready               : in  std_logic                     := 'X';             -- rready
			intel_niosv_g_0_instruction_manager_awaddr        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			intel_niosv_g_0_instruction_manager_awlen         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- awlen
			intel_niosv_g_0_instruction_manager_awsize        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			intel_niosv_g_0_instruction_manager_awburst       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			intel_niosv_g_0_instruction_manager_awprot        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			intel_niosv_g_0_instruction_manager_awvalid       : in  std_logic                     := 'X';             -- awvalid
			intel_niosv_g_0_instruction_manager_awready       : out std_logic;                                        -- awready
			intel_niosv_g_0_instruction_manager_wdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			intel_niosv_g_0_instruction_manager_wstrb         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			intel_niosv_g_0_instruction_manager_wlast         : in  std_logic                     := 'X';             -- wlast
			intel_niosv_g_0_instruction_manager_wvalid        : in  std_logic                     := 'X';             -- wvalid
			intel_niosv_g_0_instruction_manager_wready        : out std_logic;                                        -- wready
			intel_niosv_g_0_instruction_manager_bresp         : out std_logic_vector(1 downto 0);                     -- bresp
			intel_niosv_g_0_instruction_manager_bvalid        : out std_logic;                                        -- bvalid
			intel_niosv_g_0_instruction_manager_bready        : in  std_logic                     := 'X';             -- bready
			intel_niosv_g_0_instruction_manager_araddr        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			intel_niosv_g_0_instruction_manager_arlen         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- arlen
			intel_niosv_g_0_instruction_manager_arsize        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			intel_niosv_g_0_instruction_manager_arburst       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			intel_niosv_g_0_instruction_manager_arprot        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			intel_niosv_g_0_instruction_manager_arvalid       : in  std_logic                     := 'X';             -- arvalid
			intel_niosv_g_0_instruction_manager_arready       : out std_logic;                                        -- arready
			intel_niosv_g_0_instruction_manager_rdata         : out std_logic_vector(31 downto 0);                    -- rdata
			intel_niosv_g_0_instruction_manager_rresp         : out std_logic_vector(1 downto 0);                     -- rresp
			intel_niosv_g_0_instruction_manager_rlast         : out std_logic;                                        -- rlast
			intel_niosv_g_0_instruction_manager_rvalid        : out std_logic;                                        -- rvalid
			intel_niosv_g_0_instruction_manager_rready        : in  std_logic                     := 'X';             -- rready
			clk_50_out_clk_clk                                : in  std_logic                     := 'X';             -- clk
			intel_niosv_g_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			bt0_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			bt0_s1_write                                      : out std_logic;                                        -- write
			bt0_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			bt0_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			bt0_s1_chipselect                                 : out std_logic;                                        -- chipselect
			i2c_opencores_0_avalon_slave_0_address            : out std_logic_vector(2 downto 0);                     -- address
			i2c_opencores_0_avalon_slave_0_write              : out std_logic;                                        -- write
			i2c_opencores_0_avalon_slave_0_readdata           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_opencores_0_avalon_slave_0_writedata          : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_opencores_0_avalon_slave_0_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect         : out std_logic;                                        -- chipselect
			intel_niosv_g_0_dm_agent_address                  : out std_logic_vector(15 downto 0);                    -- address
			intel_niosv_g_0_dm_agent_write                    : out std_logic;                                        -- write
			intel_niosv_g_0_dm_agent_read                     : out std_logic;                                        -- read
			intel_niosv_g_0_dm_agent_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			intel_niosv_g_0_dm_agent_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			intel_niosv_g_0_dm_agent_readdatavalid            : in  std_logic                     := 'X';             -- readdatavalid
			intel_niosv_g_0_dm_agent_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			intel_niosv_g_0_timer_sw_agent_address            : out std_logic_vector(5 downto 0);                     -- address
			intel_niosv_g_0_timer_sw_agent_write              : out std_logic;                                        -- write
			intel_niosv_g_0_timer_sw_agent_read               : out std_logic;                                        -- read
			intel_niosv_g_0_timer_sw_agent_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			intel_niosv_g_0_timer_sw_agent_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			intel_niosv_g_0_timer_sw_agent_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			intel_niosv_g_0_timer_sw_agent_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			intel_niosv_g_0_timer_sw_agent_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write               : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect          : out std_logic;                                        -- chipselect
			led0_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			led0_s1_write                                     : out std_logic;                                        -- write
			led0_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led0_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			led0_s1_chipselect                                : out std_logic;                                        -- chipselect
			mm_clock_crossing_bridge_0_s0_address             : out std_logic_vector(25 downto 0);                    -- address
			mm_clock_crossing_bridge_0_s0_write               : out std_logic;                                        -- write
			mm_clock_crossing_bridge_0_s0_read                : out std_logic;                                        -- read
			mm_clock_crossing_bridge_0_s0_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mm_clock_crossing_bridge_0_s0_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			mm_clock_crossing_bridge_0_s0_burstcount          : out std_logic_vector(0 downto 0);                     -- burstcount
			mm_clock_crossing_bridge_0_s0_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_clock_crossing_bridge_0_s0_readdatavalid       : in  std_logic                     := 'X';             -- readdatavalid
			mm_clock_crossing_bridge_0_s0_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			mm_clock_crossing_bridge_0_s0_debugaccess         : out std_logic;                                        -- debugaccess
			ram_0_s1_address                                  : out std_logic_vector(14 downto 0);                    -- address
			ram_0_s1_write                                    : out std_logic;                                        -- write
			ram_0_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ram_0_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			ram_0_s1_byteenable                               : out std_logic_vector(3 downto 0);                     -- byteenable
			ram_0_s1_chipselect                               : out std_logic;                                        -- chipselect
			ram_0_s1_clken                                    : out std_logic;                                        -- clken
			rh_temp_drdy_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			rh_temp_drdy_s1_write                             : out std_logic;                                        -- write
			rh_temp_drdy_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rh_temp_drdy_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			rh_temp_drdy_s1_chipselect                        : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component NIOS_RFS2_mm_interconnect_0;

	component NIOS_RFS2_mm_interconnect_2 is
		port (
			clk_100_out_clk_clk                           : in  std_logic                     := 'X';             -- clk
			mm_bridge_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mm_bridge_0_m0_address                        : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			mm_bridge_0_m0_waitrequest                    : out std_logic;                                        -- waitrequest
			mm_bridge_0_m0_burstcount                     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			mm_bridge_0_m0_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mm_bridge_0_m0_read                           : in  std_logic                     := 'X';             -- read
			mm_bridge_0_m0_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			mm_bridge_0_m0_readdatavalid                  : out std_logic;                                        -- readdatavalid
			mm_bridge_0_m0_write                          : in  std_logic                     := 'X';             -- write
			mm_bridge_0_m0_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_bridge_0_m0_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			SDRAM_s1_address                              : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_s1_write                                : out std_logic;                                        -- write
			SDRAM_s1_read                                 : out std_logic;                                        -- read
			SDRAM_s1_readdata                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                            : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_s1_byteenable                           : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                        : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                           : out std_logic                                         -- chipselect
		);
	end component NIOS_RFS2_mm_interconnect_2;

	component NIOS_RFS2_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(15 downto 0)         -- irq
		);
	end component NIOS_RFS2_irq_mapper;

	component nios_rfs2_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_rfs2_rst_controller;

	component nios_rfs2_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_rfs2_rst_controller_001;

	signal mm_clock_crossing_bridge_0_m0_waitrequest                       : std_logic;                     -- mm_bridge_0:s0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	signal mm_clock_crossing_bridge_0_m0_readdata                          : std_logic_vector(31 downto 0); -- mm_bridge_0:s0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	signal mm_clock_crossing_bridge_0_m0_debugaccess                       : std_logic;                     -- mm_clock_crossing_bridge_0:m0_debugaccess -> mm_bridge_0:s0_debugaccess
	signal mm_clock_crossing_bridge_0_m0_address                           : std_logic_vector(25 downto 0); -- mm_clock_crossing_bridge_0:m0_address -> mm_bridge_0:s0_address
	signal mm_clock_crossing_bridge_0_m0_read                              : std_logic;                     -- mm_clock_crossing_bridge_0:m0_read -> mm_bridge_0:s0_read
	signal mm_clock_crossing_bridge_0_m0_byteenable                        : std_logic_vector(3 downto 0);  -- mm_clock_crossing_bridge_0:m0_byteenable -> mm_bridge_0:s0_byteenable
	signal mm_clock_crossing_bridge_0_m0_readdatavalid                     : std_logic;                     -- mm_bridge_0:s0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	signal mm_clock_crossing_bridge_0_m0_writedata                         : std_logic_vector(31 downto 0); -- mm_clock_crossing_bridge_0:m0_writedata -> mm_bridge_0:s0_writedata
	signal mm_clock_crossing_bridge_0_m0_write                             : std_logic;                     -- mm_clock_crossing_bridge_0:m0_write -> mm_bridge_0:s0_write
	signal mm_clock_crossing_bridge_0_m0_burstcount                        : std_logic_vector(0 downto 0);  -- mm_clock_crossing_bridge_0:m0_burstcount -> mm_bridge_0:s0_burstcount
	signal intel_niosv_g_0_data_manager_arlen                              : std_logic_vector(7 downto 0);  -- intel_niosv_g_0:data_manager_arlen -> mm_interconnect_0:intel_niosv_g_0_data_manager_arlen
	signal intel_niosv_g_0_data_manager_wstrb                              : std_logic_vector(3 downto 0);  -- intel_niosv_g_0:data_manager_wstrb -> mm_interconnect_0:intel_niosv_g_0_data_manager_wstrb
	signal intel_niosv_g_0_data_manager_wready                             : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_data_manager_wready -> intel_niosv_g_0:data_manager_wready
	signal intel_niosv_g_0_data_manager_rready                             : std_logic;                     -- intel_niosv_g_0:data_manager_rready -> mm_interconnect_0:intel_niosv_g_0_data_manager_rready
	signal intel_niosv_g_0_data_manager_awlen                              : std_logic_vector(7 downto 0);  -- intel_niosv_g_0:data_manager_awlen -> mm_interconnect_0:intel_niosv_g_0_data_manager_awlen
	signal intel_niosv_g_0_data_manager_wvalid                             : std_logic;                     -- intel_niosv_g_0:data_manager_wvalid -> mm_interconnect_0:intel_niosv_g_0_data_manager_wvalid
	signal intel_niosv_g_0_data_manager_araddr                             : std_logic_vector(31 downto 0); -- intel_niosv_g_0:data_manager_araddr -> mm_interconnect_0:intel_niosv_g_0_data_manager_araddr
	signal intel_niosv_g_0_data_manager_arprot                             : std_logic_vector(2 downto 0);  -- intel_niosv_g_0:data_manager_arprot -> mm_interconnect_0:intel_niosv_g_0_data_manager_arprot
	signal intel_niosv_g_0_data_manager_awprot                             : std_logic_vector(2 downto 0);  -- intel_niosv_g_0:data_manager_awprot -> mm_interconnect_0:intel_niosv_g_0_data_manager_awprot
	signal intel_niosv_g_0_data_manager_wdata                              : std_logic_vector(31 downto 0); -- intel_niosv_g_0:data_manager_wdata -> mm_interconnect_0:intel_niosv_g_0_data_manager_wdata
	signal intel_niosv_g_0_data_manager_arvalid                            : std_logic;                     -- intel_niosv_g_0:data_manager_arvalid -> mm_interconnect_0:intel_niosv_g_0_data_manager_arvalid
	signal intel_niosv_g_0_data_manager_awaddr                             : std_logic_vector(31 downto 0); -- intel_niosv_g_0:data_manager_awaddr -> mm_interconnect_0:intel_niosv_g_0_data_manager_awaddr
	signal intel_niosv_g_0_data_manager_bresp                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:intel_niosv_g_0_data_manager_bresp -> intel_niosv_g_0:data_manager_bresp
	signal intel_niosv_g_0_data_manager_arready                            : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_data_manager_arready -> intel_niosv_g_0:data_manager_arready
	signal intel_niosv_g_0_data_manager_rdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:intel_niosv_g_0_data_manager_rdata -> intel_niosv_g_0:data_manager_rdata
	signal intel_niosv_g_0_data_manager_awready                            : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_data_manager_awready -> intel_niosv_g_0:data_manager_awready
	signal intel_niosv_g_0_data_manager_arsize                             : std_logic_vector(2 downto 0);  -- intel_niosv_g_0:data_manager_arsize -> mm_interconnect_0:intel_niosv_g_0_data_manager_arsize
	signal intel_niosv_g_0_data_manager_rlast                              : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_data_manager_rlast -> intel_niosv_g_0:data_manager_rlast
	signal intel_niosv_g_0_data_manager_bready                             : std_logic;                     -- intel_niosv_g_0:data_manager_bready -> mm_interconnect_0:intel_niosv_g_0_data_manager_bready
	signal intel_niosv_g_0_data_manager_wlast                              : std_logic;                     -- intel_niosv_g_0:data_manager_wlast -> mm_interconnect_0:intel_niosv_g_0_data_manager_wlast
	signal intel_niosv_g_0_data_manager_rresp                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:intel_niosv_g_0_data_manager_rresp -> intel_niosv_g_0:data_manager_rresp
	signal intel_niosv_g_0_data_manager_bvalid                             : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_data_manager_bvalid -> intel_niosv_g_0:data_manager_bvalid
	signal intel_niosv_g_0_data_manager_awsize                             : std_logic_vector(2 downto 0);  -- intel_niosv_g_0:data_manager_awsize -> mm_interconnect_0:intel_niosv_g_0_data_manager_awsize
	signal intel_niosv_g_0_data_manager_awvalid                            : std_logic;                     -- intel_niosv_g_0:data_manager_awvalid -> mm_interconnect_0:intel_niosv_g_0_data_manager_awvalid
	signal intel_niosv_g_0_data_manager_rvalid                             : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_data_manager_rvalid -> intel_niosv_g_0:data_manager_rvalid
	signal intel_niosv_g_0_instruction_manager_awburst                     : std_logic_vector(1 downto 0);  -- intel_niosv_g_0:instruction_manager_awburst -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awburst
	signal intel_niosv_g_0_instruction_manager_arlen                       : std_logic_vector(7 downto 0);  -- intel_niosv_g_0:instruction_manager_arlen -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arlen
	signal intel_niosv_g_0_instruction_manager_wstrb                       : std_logic_vector(3 downto 0);  -- intel_niosv_g_0:instruction_manager_wstrb -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_wstrb
	signal intel_niosv_g_0_instruction_manager_wready                      : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_wready -> intel_niosv_g_0:instruction_manager_wready
	signal intel_niosv_g_0_instruction_manager_rready                      : std_logic;                     -- intel_niosv_g_0:instruction_manager_rready -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_rready
	signal intel_niosv_g_0_instruction_manager_awlen                       : std_logic_vector(7 downto 0);  -- intel_niosv_g_0:instruction_manager_awlen -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awlen
	signal intel_niosv_g_0_instruction_manager_wvalid                      : std_logic;                     -- intel_niosv_g_0:instruction_manager_wvalid -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_wvalid
	signal intel_niosv_g_0_instruction_manager_araddr                      : std_logic_vector(31 downto 0); -- intel_niosv_g_0:instruction_manager_araddr -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_araddr
	signal intel_niosv_g_0_instruction_manager_arprot                      : std_logic_vector(2 downto 0);  -- intel_niosv_g_0:instruction_manager_arprot -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arprot
	signal intel_niosv_g_0_instruction_manager_awprot                      : std_logic_vector(2 downto 0);  -- intel_niosv_g_0:instruction_manager_awprot -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awprot
	signal intel_niosv_g_0_instruction_manager_wdata                       : std_logic_vector(31 downto 0); -- intel_niosv_g_0:instruction_manager_wdata -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_wdata
	signal intel_niosv_g_0_instruction_manager_arvalid                     : std_logic;                     -- intel_niosv_g_0:instruction_manager_arvalid -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arvalid
	signal intel_niosv_g_0_instruction_manager_awaddr                      : std_logic_vector(31 downto 0); -- intel_niosv_g_0:instruction_manager_awaddr -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awaddr
	signal intel_niosv_g_0_instruction_manager_bresp                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_bresp -> intel_niosv_g_0:instruction_manager_bresp
	signal intel_niosv_g_0_instruction_manager_arready                     : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_arready -> intel_niosv_g_0:instruction_manager_arready
	signal intel_niosv_g_0_instruction_manager_rdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_rdata -> intel_niosv_g_0:instruction_manager_rdata
	signal intel_niosv_g_0_instruction_manager_arburst                     : std_logic_vector(1 downto 0);  -- intel_niosv_g_0:instruction_manager_arburst -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arburst
	signal intel_niosv_g_0_instruction_manager_awready                     : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_awready -> intel_niosv_g_0:instruction_manager_awready
	signal intel_niosv_g_0_instruction_manager_arsize                      : std_logic_vector(2 downto 0);  -- intel_niosv_g_0:instruction_manager_arsize -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arsize
	signal intel_niosv_g_0_instruction_manager_rlast                       : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_rlast -> intel_niosv_g_0:instruction_manager_rlast
	signal intel_niosv_g_0_instruction_manager_bready                      : std_logic;                     -- intel_niosv_g_0:instruction_manager_bready -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_bready
	signal intel_niosv_g_0_instruction_manager_wlast                       : std_logic;                     -- intel_niosv_g_0:instruction_manager_wlast -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_wlast
	signal intel_niosv_g_0_instruction_manager_rresp                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_rresp -> intel_niosv_g_0:instruction_manager_rresp
	signal intel_niosv_g_0_instruction_manager_bvalid                      : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_bvalid -> intel_niosv_g_0:instruction_manager_bvalid
	signal intel_niosv_g_0_instruction_manager_awsize                      : std_logic_vector(2 downto 0);  -- intel_niosv_g_0:instruction_manager_awsize -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awsize
	signal intel_niosv_g_0_instruction_manager_awvalid                     : std_logic;                     -- intel_niosv_g_0:instruction_manager_awvalid -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awvalid
	signal intel_niosv_g_0_instruction_manager_rvalid                      : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_instruction_manager_rvalid -> intel_niosv_g_0:instruction_manager_rvalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect     : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata       : std_logic_vector(7 downto 0);  -- i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	signal i2c_opencores_0_avalon_slave_0_waitrequest                      : std_logic;                     -- i2c_opencores_0:wb_ack_o -> i2c_opencores_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata      : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_intel_niosv_g_0_dm_agent_readdata             : std_logic_vector(31 downto 0); -- intel_niosv_g_0:dm_agent_readdata -> mm_interconnect_0:intel_niosv_g_0_dm_agent_readdata
	signal mm_interconnect_0_intel_niosv_g_0_dm_agent_waitrequest          : std_logic;                     -- intel_niosv_g_0:dm_agent_waitrequest -> mm_interconnect_0:intel_niosv_g_0_dm_agent_waitrequest
	signal mm_interconnect_0_intel_niosv_g_0_dm_agent_address              : std_logic_vector(15 downto 0); -- mm_interconnect_0:intel_niosv_g_0_dm_agent_address -> intel_niosv_g_0:dm_agent_address
	signal mm_interconnect_0_intel_niosv_g_0_dm_agent_read                 : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_dm_agent_read -> intel_niosv_g_0:dm_agent_read
	signal mm_interconnect_0_intel_niosv_g_0_dm_agent_readdatavalid        : std_logic;                     -- intel_niosv_g_0:dm_agent_readdatavalid -> mm_interconnect_0:intel_niosv_g_0_dm_agent_readdatavalid
	signal mm_interconnect_0_intel_niosv_g_0_dm_agent_write                : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_dm_agent_write -> intel_niosv_g_0:dm_agent_write
	signal mm_interconnect_0_intel_niosv_g_0_dm_agent_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:intel_niosv_g_0_dm_agent_writedata -> intel_niosv_g_0:dm_agent_writedata
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata        : std_logic_vector(31 downto 0); -- mm_clock_crossing_bridge_0:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdata
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest     : std_logic;                     -- mm_clock_crossing_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_waitrequest
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess     : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address         : std_logic_vector(25 downto 0); -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_address -> mm_clock_crossing_bridge_0:s0_address
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read            : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_read -> mm_clock_crossing_bridge_0:s0_read
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid   : std_logic;                     -- mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdatavalid
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write           : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_write -> mm_clock_crossing_bridge_0:s0_write
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	signal mm_interconnect_0_ram_0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:ram_0_s1_chipselect -> ram_0:chipselect
	signal mm_interconnect_0_ram_0_s1_readdata                             : std_logic_vector(31 downto 0); -- ram_0:readdata -> mm_interconnect_0:ram_0_s1_readdata
	signal mm_interconnect_0_ram_0_s1_address                              : std_logic_vector(14 downto 0); -- mm_interconnect_0:ram_0_s1_address -> ram_0:address
	signal mm_interconnect_0_ram_0_s1_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ram_0_s1_byteenable -> ram_0:byteenable
	signal mm_interconnect_0_ram_0_s1_write                                : std_logic;                     -- mm_interconnect_0:ram_0_s1_write -> ram_0:write
	signal mm_interconnect_0_ram_0_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:ram_0_s1_writedata -> ram_0:writedata
	signal mm_interconnect_0_ram_0_s1_clken                                : std_logic;                     -- mm_interconnect_0:ram_0_s1_clken -> ram_0:clken
	signal mm_interconnect_0_led0_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:led0_s1_chipselect -> led0:chipselect
	signal mm_interconnect_0_led0_s1_readdata                              : std_logic_vector(31 downto 0); -- led0:readdata -> mm_interconnect_0:led0_s1_readdata
	signal mm_interconnect_0_led0_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led0_s1_address -> led0:address
	signal mm_interconnect_0_led0_s1_write                                 : std_logic;                     -- mm_interconnect_0:led0_s1_write -> mm_interconnect_0_led0_s1_write:in
	signal mm_interconnect_0_led0_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:led0_s1_writedata -> led0:writedata
	signal mm_interconnect_0_bt0_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:bt0_s1_chipselect -> bt0:chipselect
	signal mm_interconnect_0_bt0_s1_readdata                               : std_logic_vector(31 downto 0); -- bt0:readdata -> mm_interconnect_0:bt0_s1_readdata
	signal mm_interconnect_0_bt0_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:bt0_s1_address -> bt0:address
	signal mm_interconnect_0_bt0_s1_write                                  : std_logic;                     -- mm_interconnect_0:bt0_s1_write -> mm_interconnect_0_bt0_s1_write:in
	signal mm_interconnect_0_bt0_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:bt0_s1_writedata -> bt0:writedata
	signal mm_interconnect_0_rh_temp_drdy_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:rh_temp_drdy_s1_chipselect -> rh_temp_drdy:chipselect
	signal mm_interconnect_0_rh_temp_drdy_s1_readdata                      : std_logic_vector(31 downto 0); -- rh_temp_drdy:readdata -> mm_interconnect_0:rh_temp_drdy_s1_readdata
	signal mm_interconnect_0_rh_temp_drdy_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:rh_temp_drdy_s1_address -> rh_temp_drdy:address
	signal mm_interconnect_0_rh_temp_drdy_s1_write                         : std_logic;                     -- mm_interconnect_0:rh_temp_drdy_s1_write -> mm_interconnect_0_rh_temp_drdy_s1_write:in
	signal mm_interconnect_0_rh_temp_drdy_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:rh_temp_drdy_s1_writedata -> rh_temp_drdy:writedata
	signal mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdata       : std_logic_vector(31 downto 0); -- intel_niosv_g_0:timer_sw_agent_readdata -> mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_readdata
	signal mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_waitrequest    : std_logic;                     -- intel_niosv_g_0:timer_sw_agent_waitrequest -> mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_waitrequest
	signal mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_address        : std_logic_vector(5 downto 0);  -- mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_address -> intel_niosv_g_0:timer_sw_agent_address
	signal mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_read           : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_read -> intel_niosv_g_0:timer_sw_agent_read
	signal mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_byteenable     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_byteenable -> intel_niosv_g_0:timer_sw_agent_byteenable
	signal mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdatavalid  : std_logic;                     -- intel_niosv_g_0:timer_sw_agent_readdatavalid -> mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_readdatavalid
	signal mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_write          : std_logic;                     -- mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_write -> intel_niosv_g_0:timer_sw_agent_write
	signal mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_writedata -> intel_niosv_g_0:timer_sw_agent_writedata
	signal mm_bridge_0_m0_waitrequest                                      : std_logic;                     -- mm_interconnect_2:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	signal mm_bridge_0_m0_readdata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_2:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	signal mm_bridge_0_m0_debugaccess                                      : std_logic;                     -- mm_bridge_0:m0_debugaccess -> mm_interconnect_2:mm_bridge_0_m0_debugaccess
	signal mm_bridge_0_m0_address                                          : std_logic_vector(25 downto 0); -- mm_bridge_0:m0_address -> mm_interconnect_2:mm_bridge_0_m0_address
	signal mm_bridge_0_m0_read                                             : std_logic;                     -- mm_bridge_0:m0_read -> mm_interconnect_2:mm_bridge_0_m0_read
	signal mm_bridge_0_m0_byteenable                                       : std_logic_vector(3 downto 0);  -- mm_bridge_0:m0_byteenable -> mm_interconnect_2:mm_bridge_0_m0_byteenable
	signal mm_bridge_0_m0_readdatavalid                                    : std_logic;                     -- mm_interconnect_2:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	signal mm_bridge_0_m0_writedata                                        : std_logic_vector(31 downto 0); -- mm_bridge_0:m0_writedata -> mm_interconnect_2:mm_bridge_0_m0_writedata
	signal mm_bridge_0_m0_write                                            : std_logic;                     -- mm_bridge_0:m0_write -> mm_interconnect_2:mm_bridge_0_m0_write
	signal mm_bridge_0_m0_burstcount                                       : std_logic_vector(0 downto 0);  -- mm_bridge_0:m0_burstcount -> mm_interconnect_2:mm_bridge_0_m0_burstcount
	signal mm_interconnect_2_sdram_s1_chipselect                           : std_logic;                     -- mm_interconnect_2:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_2_sdram_s1_readdata                             : std_logic_vector(15 downto 0); -- SDRAM:za_data -> mm_interconnect_2:SDRAM_s1_readdata
	signal mm_interconnect_2_sdram_s1_waitrequest                          : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_2:SDRAM_s1_waitrequest
	signal mm_interconnect_2_sdram_s1_address                              : std_logic_vector(24 downto 0); -- mm_interconnect_2:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_2_sdram_s1_read                                 : std_logic;                     -- mm_interconnect_2:SDRAM_s1_read -> mm_interconnect_2_sdram_s1_read:in
	signal mm_interconnect_2_sdram_s1_byteenable                           : std_logic_vector(1 downto 0);  -- mm_interconnect_2:SDRAM_s1_byteenable -> mm_interconnect_2_sdram_s1_byteenable:in
	signal mm_interconnect_2_sdram_s1_readdatavalid                        : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_2:SDRAM_s1_readdatavalid
	signal mm_interconnect_2_sdram_s1_write                                : std_logic;                     -- mm_interconnect_2:SDRAM_s1_write -> mm_interconnect_2_sdram_s1_write:in
	signal mm_interconnect_2_sdram_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_2:SDRAM_s1_writedata -> SDRAM:az_data
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- i2c_opencores_0:wb_inta_o -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- bt0:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- rh_temp_drdy:irq -> irq_mapper:receiver3_irq
	signal intel_niosv_g_0_platform_irq_rx_irq                             : std_logic_vector(15 downto 0); -- irq_mapper:sender_irq -> intel_niosv_g_0:platform_irq_rx_irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [i2c_opencores_0:wb_rst_i, intel_niosv_g_0:ndm_reset_in_reset, intel_niosv_g_0:reset_reset, irq_mapper:reset, mm_clock_crossing_bridge_0:s0_reset, mm_interconnect_0:intel_niosv_g_0_reset_reset_bridge_in_reset_reset, ram_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [ram_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal intel_niosv_g_0_dbg_reset_out_reset                             : std_logic;                     -- intel_niosv_g_0:dbg_reset_out_reset -> rst_controller_001:reset_in0
	signal reset_bridge_100_in_reset_reset_n_ports_inv                     : std_logic;                     -- reset_bridge_100_in_reset_reset_n:inv -> [mm_bridge_0:reset, mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_2:mm_bridge_0_reset_reset_bridge_in_reset_reset]
	signal reset_bridge_50_in_reset_reset_n_ports_inv                      : std_logic;                     -- reset_bridge_50_in_reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in1]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv            : std_logic;                     -- i2c_opencores_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_led0_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_led0_s1_write:inv -> led0:write_n
	signal mm_interconnect_0_bt0_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_bt0_s1_write:inv -> bt0:write_n
	signal mm_interconnect_0_rh_temp_drdy_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_rh_temp_drdy_s1_write:inv -> rh_temp_drdy:write_n
	signal mm_interconnect_2_sdram_s1_read_ports_inv                       : std_logic;                     -- mm_interconnect_2_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_2_sdram_s1_byteenable_ports_inv                 : std_logic_vector(1 downto 0);  -- mm_interconnect_2_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_2_sdram_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_2_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [bt0:reset_n, led0:reset_n, rh_temp_drdy:reset_n, sysid_qsys_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> jtag_uart_0:rst_n

begin

	sdram : component NIOS_RFS2_SDRAM
		port map (
			clk            => clk_100_in_clk_clk,                              --                 clk.clk
			reset_n        => reset_bridge_100_in_reset_reset_n,               --               reset.reset_n
			az_addr        => mm_interconnect_2_sdram_s1_address,              --                  s1.address
			az_be_n        => mm_interconnect_2_sdram_s1_byteenable_ports_inv, --                    .byteenable_n
			az_cs          => mm_interconnect_2_sdram_s1_chipselect,           --                    .chipselect
			az_data        => mm_interconnect_2_sdram_s1_writedata,            --                    .writedata
			az_rd_n        => mm_interconnect_2_sdram_s1_read_ports_inv,       --                    .read_n
			az_wr_n        => mm_interconnect_2_sdram_s1_write_ports_inv,      --                    .write_n
			za_data        => mm_interconnect_2_sdram_s1_readdata,             --                    .readdata
			za_valid       => mm_interconnect_2_sdram_s1_readdatavalid,        --                    .readdatavalid
			za_waitrequest => mm_interconnect_2_sdram_s1_waitrequest,          --                    .waitrequest
			zs_addr        => sdram_addr,                                      -- external_connection.export
			zs_ba          => sdram_ba,                                        --                    .export
			zs_cas_n       => sdram_cas_n,                                     --                    .export
			zs_cke         => sdram_cke,                                       --                    .export
			zs_cs_n        => sdram_cs_n,                                      --                    .export
			zs_dq          => sdram_dq,                                        --                    .export
			zs_dqm         => sdram_dqm,                                       --                    .export
			zs_ras_n       => sdram_ras_n,                                     --                    .export
			zs_we_n        => sdram_we_n                                       --                    .export
		);

	bt0 : component NIOS_RFS2_bt0
		port map (
			clk        => clk_50_in_clk_clk,                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_bt0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_bt0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_bt0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_bt0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_bt0_s1_readdata,        --                    .readdata
			in_port    => bt0_export,                               -- external_connection.export
			irq        => irq_mapper_receiver2_irq                  --                 irq.irq
		);

	i2c_opencores_0 : component i2c_opencores
		port map (
			wb_clk_i   => clk_50_in_clk_clk,                                           --            clock.clk
			wb_rst_i   => rst_controller_reset_out_reset,                              --      clock_reset.reset
			scl_pad_io => i2c_scl_pad_io,                                              --           export.export
			sda_pad_io => i2c_sda_pad_io,                                              --                 .export
			wb_adr_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_opencores_0_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			wb_inta_o  => irq_mapper_receiver0_irq                                     -- interrupt_sender.irq
		);

	intel_niosv_g_0 : component NIOS_RFS2_intel_niosv_g_0
		port map (
			clk                          => clk_50_in_clk_clk,                                              --                 clk.clk
			reset_reset                  => rst_controller_reset_out_reset,                                 --               reset.reset
			instruction_manager_awsize   => intel_niosv_g_0_instruction_manager_awsize,                     -- instruction_manager.awsize
			instruction_manager_awlen    => intel_niosv_g_0_instruction_manager_awlen,                      --                    .awlen
			instruction_manager_awburst  => intel_niosv_g_0_instruction_manager_awburst,                    --                    .awburst
			instruction_manager_wlast    => intel_niosv_g_0_instruction_manager_wlast,                      --                    .wlast
			instruction_manager_arsize   => intel_niosv_g_0_instruction_manager_arsize,                     --                    .arsize
			instruction_manager_arlen    => intel_niosv_g_0_instruction_manager_arlen,                      --                    .arlen
			instruction_manager_arburst  => intel_niosv_g_0_instruction_manager_arburst,                    --                    .arburst
			instruction_manager_rlast    => intel_niosv_g_0_instruction_manager_rlast,                      --                    .rlast
			instruction_manager_awaddr   => intel_niosv_g_0_instruction_manager_awaddr,                     --                    .awaddr
			instruction_manager_awprot   => intel_niosv_g_0_instruction_manager_awprot,                     --                    .awprot
			instruction_manager_awvalid  => intel_niosv_g_0_instruction_manager_awvalid,                    --                    .awvalid
			instruction_manager_awready  => intel_niosv_g_0_instruction_manager_awready,                    --                    .awready
			instruction_manager_wdata    => intel_niosv_g_0_instruction_manager_wdata,                      --                    .wdata
			instruction_manager_wstrb    => intel_niosv_g_0_instruction_manager_wstrb,                      --                    .wstrb
			instruction_manager_wvalid   => intel_niosv_g_0_instruction_manager_wvalid,                     --                    .wvalid
			instruction_manager_wready   => intel_niosv_g_0_instruction_manager_wready,                     --                    .wready
			instruction_manager_bresp    => intel_niosv_g_0_instruction_manager_bresp,                      --                    .bresp
			instruction_manager_bvalid   => intel_niosv_g_0_instruction_manager_bvalid,                     --                    .bvalid
			instruction_manager_bready   => intel_niosv_g_0_instruction_manager_bready,                     --                    .bready
			instruction_manager_araddr   => intel_niosv_g_0_instruction_manager_araddr,                     --                    .araddr
			instruction_manager_arprot   => intel_niosv_g_0_instruction_manager_arprot,                     --                    .arprot
			instruction_manager_arvalid  => intel_niosv_g_0_instruction_manager_arvalid,                    --                    .arvalid
			instruction_manager_arready  => intel_niosv_g_0_instruction_manager_arready,                    --                    .arready
			instruction_manager_rdata    => intel_niosv_g_0_instruction_manager_rdata,                      --                    .rdata
			instruction_manager_rresp    => intel_niosv_g_0_instruction_manager_rresp,                      --                    .rresp
			instruction_manager_rvalid   => intel_niosv_g_0_instruction_manager_rvalid,                     --                    .rvalid
			instruction_manager_rready   => intel_niosv_g_0_instruction_manager_rready,                     --                    .rready
			data_manager_awsize          => intel_niosv_g_0_data_manager_awsize,                            --        data_manager.awsize
			data_manager_awlen           => intel_niosv_g_0_data_manager_awlen,                             --                    .awlen
			data_manager_wlast           => intel_niosv_g_0_data_manager_wlast,                             --                    .wlast
			data_manager_arsize          => intel_niosv_g_0_data_manager_arsize,                            --                    .arsize
			data_manager_arlen           => intel_niosv_g_0_data_manager_arlen,                             --                    .arlen
			data_manager_rlast           => intel_niosv_g_0_data_manager_rlast,                             --                    .rlast
			data_manager_awaddr          => intel_niosv_g_0_data_manager_awaddr,                            --                    .awaddr
			data_manager_awprot          => intel_niosv_g_0_data_manager_awprot,                            --                    .awprot
			data_manager_awvalid         => intel_niosv_g_0_data_manager_awvalid,                           --                    .awvalid
			data_manager_awready         => intel_niosv_g_0_data_manager_awready,                           --                    .awready
			data_manager_wdata           => intel_niosv_g_0_data_manager_wdata,                             --                    .wdata
			data_manager_wstrb           => intel_niosv_g_0_data_manager_wstrb,                             --                    .wstrb
			data_manager_wvalid          => intel_niosv_g_0_data_manager_wvalid,                            --                    .wvalid
			data_manager_wready          => intel_niosv_g_0_data_manager_wready,                            --                    .wready
			data_manager_bresp           => intel_niosv_g_0_data_manager_bresp,                             --                    .bresp
			data_manager_bvalid          => intel_niosv_g_0_data_manager_bvalid,                            --                    .bvalid
			data_manager_bready          => intel_niosv_g_0_data_manager_bready,                            --                    .bready
			data_manager_araddr          => intel_niosv_g_0_data_manager_araddr,                            --                    .araddr
			data_manager_arprot          => intel_niosv_g_0_data_manager_arprot,                            --                    .arprot
			data_manager_arvalid         => intel_niosv_g_0_data_manager_arvalid,                           --                    .arvalid
			data_manager_arready         => intel_niosv_g_0_data_manager_arready,                           --                    .arready
			data_manager_rdata           => intel_niosv_g_0_data_manager_rdata,                             --                    .rdata
			data_manager_rresp           => intel_niosv_g_0_data_manager_rresp,                             --                    .rresp
			data_manager_rvalid          => intel_niosv_g_0_data_manager_rvalid,                            --                    .rvalid
			data_manager_rready          => intel_niosv_g_0_data_manager_rready,                            --                    .rready
			platform_irq_rx_irq          => intel_niosv_g_0_platform_irq_rx_irq,                            --     platform_irq_rx.irq
			ndm_reset_in_reset           => rst_controller_reset_out_reset,                                 --        ndm_reset_in.reset
			timer_sw_agent_address       => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_address,       --      timer_sw_agent.address
			timer_sw_agent_byteenable    => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_byteenable,    --                    .byteenable
			timer_sw_agent_read          => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_read,          --                    .read
			timer_sw_agent_readdata      => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdata,      --                    .readdata
			timer_sw_agent_write         => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_write,         --                    .write
			timer_sw_agent_writedata     => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_writedata,     --                    .writedata
			timer_sw_agent_waitrequest   => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_waitrequest,   --                    .waitrequest
			timer_sw_agent_readdatavalid => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdatavalid, --                    .readdatavalid
			dm_agent_address             => mm_interconnect_0_intel_niosv_g_0_dm_agent_address,             --            dm_agent.address
			dm_agent_read                => mm_interconnect_0_intel_niosv_g_0_dm_agent_read,                --                    .read
			dm_agent_readdata            => mm_interconnect_0_intel_niosv_g_0_dm_agent_readdata,            --                    .readdata
			dm_agent_write               => mm_interconnect_0_intel_niosv_g_0_dm_agent_write,               --                    .write
			dm_agent_writedata           => mm_interconnect_0_intel_niosv_g_0_dm_agent_writedata,           --                    .writedata
			dm_agent_waitrequest         => mm_interconnect_0_intel_niosv_g_0_dm_agent_waitrequest,         --                    .waitrequest
			dm_agent_readdatavalid       => mm_interconnect_0_intel_niosv_g_0_dm_agent_readdatavalid,       --                    .readdatavalid
			dbg_reset_out_reset          => intel_niosv_g_0_dbg_reset_out_reset                             --       dbg_reset_out.reset
		);

	jtag_uart_0 : component altera_avalon_jtag_uart
		generic map (
			readBufferDepth            => 64,
			readIRQThreshold           => 8,
			useRegistersForReadBuffer  => false,
			useRegistersForWriteBuffer => false,
			writeBufferDepth           => 64,
			writeIRQThreshold          => 8,
			printingMethod             => false,
			FIFO_WIDTH                 => 8,
			WR_WIDTHU                  => 6,
			RD_WIDTHU                  => 6,
			write_le                   => "ON",
			read_le                    => "ON",
			HEX_WRITE_DEPTH_STR        => 64,
			HEX_READ_DEPTH_STR         => 64,
			legacySignalAllow          => false
		)
		port map (
			clk            => clk_50_in_clk_clk,                                               --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                         --               irq.irq
		);

	led0 : component NIOS_RFS2_led0
		port map (
			clk        => clk_50_in_clk_clk,                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_led0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led0_s1_readdata,        --                    .readdata
			out_port   => led_nios_export                            -- external_connection.export
		);

	mm_bridge_0 : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 26,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => clk_100_in_clk_clk,                          --   clk.clk
			reset            => reset_bridge_100_in_reset_reset_n_ports_inv, -- reset.reset
			s0_waitrequest   => mm_clock_crossing_bridge_0_m0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_clock_crossing_bridge_0_m0_readdata,      --      .readdata
			s0_readdatavalid => mm_clock_crossing_bridge_0_m0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_clock_crossing_bridge_0_m0_burstcount,    --      .burstcount
			s0_writedata     => mm_clock_crossing_bridge_0_m0_writedata,     --      .writedata
			s0_address       => mm_clock_crossing_bridge_0_m0_address,       --      .address
			s0_write         => mm_clock_crossing_bridge_0_m0_write,         --      .write
			s0_read          => mm_clock_crossing_bridge_0_m0_read,          --      .read
			s0_byteenable    => mm_clock_crossing_bridge_0_m0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_clock_crossing_bridge_0_m0_debugaccess,   --      .debugaccess
			m0_waitrequest   => mm_bridge_0_m0_waitrequest,                  --    m0.waitrequest
			m0_readdata      => mm_bridge_0_m0_readdata,                     --      .readdata
			m0_readdatavalid => mm_bridge_0_m0_readdatavalid,                --      .readdatavalid
			m0_burstcount    => mm_bridge_0_m0_burstcount,                   --      .burstcount
			m0_writedata     => mm_bridge_0_m0_writedata,                    --      .writedata
			m0_address       => mm_bridge_0_m0_address,                      --      .address
			m0_write         => mm_bridge_0_m0_write,                        --      .write
			m0_read          => mm_bridge_0_m0_read,                         --      .read
			m0_byteenable    => mm_bridge_0_m0_byteenable,                   --      .byteenable
			m0_debugaccess   => mm_bridge_0_m0_debugaccess,                  --      .debugaccess
			s0_response      => open,                                        -- (terminated)
			m0_response      => "00"                                         -- (terminated)
		);

	mm_clock_crossing_bridge_0 : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 26,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 64,
			RESPONSE_FIFO_DEPTH => 64,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => clk_100_in_clk_clk,                                            --   m0_clk.clk
			m0_reset         => reset_bridge_100_in_reset_reset_n_ports_inv,                   -- m0_reset.reset
			s0_clk           => clk_50_in_clk_clk,                                             --   s0_clk.clk
			s0_reset         => rst_controller_reset_out_reset,                                -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address,       --         .address
			s0_write         => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write,         --         .write
			s0_read          => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => mm_clock_crossing_bridge_0_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => mm_clock_crossing_bridge_0_m0_readdata,                        --         .readdata
			m0_readdatavalid => mm_clock_crossing_bridge_0_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => mm_clock_crossing_bridge_0_m0_burstcount,                      --         .burstcount
			m0_writedata     => mm_clock_crossing_bridge_0_m0_writedata,                       --         .writedata
			m0_address       => mm_clock_crossing_bridge_0_m0_address,                         --         .address
			m0_write         => mm_clock_crossing_bridge_0_m0_write,                           --         .write
			m0_read          => mm_clock_crossing_bridge_0_m0_read,                            --         .read
			m0_byteenable    => mm_clock_crossing_bridge_0_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => mm_clock_crossing_bridge_0_m0_debugaccess                      --         .debugaccess
		);

	ram_0 : component NIOS_RFS2_ram_0
		port map (
			clk        => clk_50_in_clk_clk,                     --   clk1.clk
			address    => mm_interconnect_0_ram_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,        -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,    --       .reset_req
			freeze     => '0'                                    -- (terminated)
		);

	rh_temp_drdy : component NIOS_RFS2_bt0
		port map (
			clk        => clk_50_in_clk_clk,                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_rh_temp_drdy_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_rh_temp_drdy_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_rh_temp_drdy_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_rh_temp_drdy_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_rh_temp_drdy_s1_readdata,        --                    .readdata
			in_port    => rh_temp_drdy_export,                               -- external_connection.export
			irq        => irq_mapper_receiver3_irq                           --                 irq.irq
		);

	sysid_qsys_0 : component NIOS_RFS2_sysid_qsys_0
		port map (
			clock    => clk_50_in_clk_clk,                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component NIOS_RFS2_mm_interconnect_0
		port map (
			intel_niosv_g_0_data_manager_awaddr               => intel_niosv_g_0_data_manager_awaddr,                            --                intel_niosv_g_0_data_manager.awaddr
			intel_niosv_g_0_data_manager_awlen                => intel_niosv_g_0_data_manager_awlen,                             --                                            .awlen
			intel_niosv_g_0_data_manager_awsize               => intel_niosv_g_0_data_manager_awsize,                            --                                            .awsize
			intel_niosv_g_0_data_manager_awprot               => intel_niosv_g_0_data_manager_awprot,                            --                                            .awprot
			intel_niosv_g_0_data_manager_awvalid              => intel_niosv_g_0_data_manager_awvalid,                           --                                            .awvalid
			intel_niosv_g_0_data_manager_awready              => intel_niosv_g_0_data_manager_awready,                           --                                            .awready
			intel_niosv_g_0_data_manager_wdata                => intel_niosv_g_0_data_manager_wdata,                             --                                            .wdata
			intel_niosv_g_0_data_manager_wstrb                => intel_niosv_g_0_data_manager_wstrb,                             --                                            .wstrb
			intel_niosv_g_0_data_manager_wlast                => intel_niosv_g_0_data_manager_wlast,                             --                                            .wlast
			intel_niosv_g_0_data_manager_wvalid               => intel_niosv_g_0_data_manager_wvalid,                            --                                            .wvalid
			intel_niosv_g_0_data_manager_wready               => intel_niosv_g_0_data_manager_wready,                            --                                            .wready
			intel_niosv_g_0_data_manager_bresp                => intel_niosv_g_0_data_manager_bresp,                             --                                            .bresp
			intel_niosv_g_0_data_manager_bvalid               => intel_niosv_g_0_data_manager_bvalid,                            --                                            .bvalid
			intel_niosv_g_0_data_manager_bready               => intel_niosv_g_0_data_manager_bready,                            --                                            .bready
			intel_niosv_g_0_data_manager_araddr               => intel_niosv_g_0_data_manager_araddr,                            --                                            .araddr
			intel_niosv_g_0_data_manager_arlen                => intel_niosv_g_0_data_manager_arlen,                             --                                            .arlen
			intel_niosv_g_0_data_manager_arsize               => intel_niosv_g_0_data_manager_arsize,                            --                                            .arsize
			intel_niosv_g_0_data_manager_arprot               => intel_niosv_g_0_data_manager_arprot,                            --                                            .arprot
			intel_niosv_g_0_data_manager_arvalid              => intel_niosv_g_0_data_manager_arvalid,                           --                                            .arvalid
			intel_niosv_g_0_data_manager_arready              => intel_niosv_g_0_data_manager_arready,                           --                                            .arready
			intel_niosv_g_0_data_manager_rdata                => intel_niosv_g_0_data_manager_rdata,                             --                                            .rdata
			intel_niosv_g_0_data_manager_rresp                => intel_niosv_g_0_data_manager_rresp,                             --                                            .rresp
			intel_niosv_g_0_data_manager_rlast                => intel_niosv_g_0_data_manager_rlast,                             --                                            .rlast
			intel_niosv_g_0_data_manager_rvalid               => intel_niosv_g_0_data_manager_rvalid,                            --                                            .rvalid
			intel_niosv_g_0_data_manager_rready               => intel_niosv_g_0_data_manager_rready,                            --                                            .rready
			intel_niosv_g_0_instruction_manager_awaddr        => intel_niosv_g_0_instruction_manager_awaddr,                     --         intel_niosv_g_0_instruction_manager.awaddr
			intel_niosv_g_0_instruction_manager_awlen         => intel_niosv_g_0_instruction_manager_awlen,                      --                                            .awlen
			intel_niosv_g_0_instruction_manager_awsize        => intel_niosv_g_0_instruction_manager_awsize,                     --                                            .awsize
			intel_niosv_g_0_instruction_manager_awburst       => intel_niosv_g_0_instruction_manager_awburst,                    --                                            .awburst
			intel_niosv_g_0_instruction_manager_awprot        => intel_niosv_g_0_instruction_manager_awprot,                     --                                            .awprot
			intel_niosv_g_0_instruction_manager_awvalid       => intel_niosv_g_0_instruction_manager_awvalid,                    --                                            .awvalid
			intel_niosv_g_0_instruction_manager_awready       => intel_niosv_g_0_instruction_manager_awready,                    --                                            .awready
			intel_niosv_g_0_instruction_manager_wdata         => intel_niosv_g_0_instruction_manager_wdata,                      --                                            .wdata
			intel_niosv_g_0_instruction_manager_wstrb         => intel_niosv_g_0_instruction_manager_wstrb,                      --                                            .wstrb
			intel_niosv_g_0_instruction_manager_wlast         => intel_niosv_g_0_instruction_manager_wlast,                      --                                            .wlast
			intel_niosv_g_0_instruction_manager_wvalid        => intel_niosv_g_0_instruction_manager_wvalid,                     --                                            .wvalid
			intel_niosv_g_0_instruction_manager_wready        => intel_niosv_g_0_instruction_manager_wready,                     --                                            .wready
			intel_niosv_g_0_instruction_manager_bresp         => intel_niosv_g_0_instruction_manager_bresp,                      --                                            .bresp
			intel_niosv_g_0_instruction_manager_bvalid        => intel_niosv_g_0_instruction_manager_bvalid,                     --                                            .bvalid
			intel_niosv_g_0_instruction_manager_bready        => intel_niosv_g_0_instruction_manager_bready,                     --                                            .bready
			intel_niosv_g_0_instruction_manager_araddr        => intel_niosv_g_0_instruction_manager_araddr,                     --                                            .araddr
			intel_niosv_g_0_instruction_manager_arlen         => intel_niosv_g_0_instruction_manager_arlen,                      --                                            .arlen
			intel_niosv_g_0_instruction_manager_arsize        => intel_niosv_g_0_instruction_manager_arsize,                     --                                            .arsize
			intel_niosv_g_0_instruction_manager_arburst       => intel_niosv_g_0_instruction_manager_arburst,                    --                                            .arburst
			intel_niosv_g_0_instruction_manager_arprot        => intel_niosv_g_0_instruction_manager_arprot,                     --                                            .arprot
			intel_niosv_g_0_instruction_manager_arvalid       => intel_niosv_g_0_instruction_manager_arvalid,                    --                                            .arvalid
			intel_niosv_g_0_instruction_manager_arready       => intel_niosv_g_0_instruction_manager_arready,                    --                                            .arready
			intel_niosv_g_0_instruction_manager_rdata         => intel_niosv_g_0_instruction_manager_rdata,                      --                                            .rdata
			intel_niosv_g_0_instruction_manager_rresp         => intel_niosv_g_0_instruction_manager_rresp,                      --                                            .rresp
			intel_niosv_g_0_instruction_manager_rlast         => intel_niosv_g_0_instruction_manager_rlast,                      --                                            .rlast
			intel_niosv_g_0_instruction_manager_rvalid        => intel_niosv_g_0_instruction_manager_rvalid,                     --                                            .rvalid
			intel_niosv_g_0_instruction_manager_rready        => intel_niosv_g_0_instruction_manager_rready,                     --                                            .rready
			clk_50_out_clk_clk                                => clk_50_in_clk_clk,                                              --                              clk_50_out_clk.clk
			intel_niosv_g_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                 -- intel_niosv_g_0_reset_reset_bridge_in_reset.reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset     => rst_controller_001_reset_out_reset,                             --     jtag_uart_0_reset_reset_bridge_in_reset.reset
			bt0_s1_address                                    => mm_interconnect_0_bt0_s1_address,                               --                                      bt0_s1.address
			bt0_s1_write                                      => mm_interconnect_0_bt0_s1_write,                                 --                                            .write
			bt0_s1_readdata                                   => mm_interconnect_0_bt0_s1_readdata,                              --                                            .readdata
			bt0_s1_writedata                                  => mm_interconnect_0_bt0_s1_writedata,                             --                                            .writedata
			bt0_s1_chipselect                                 => mm_interconnect_0_bt0_s1_chipselect,                            --                                            .chipselect
			i2c_opencores_0_avalon_slave_0_address            => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,       --              i2c_opencores_0_avalon_slave_0.address
			i2c_opencores_0_avalon_slave_0_write              => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,         --                                            .write
			i2c_opencores_0_avalon_slave_0_readdata           => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,      --                                            .readdata
			i2c_opencores_0_avalon_slave_0_writedata          => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,     --                                            .writedata
			i2c_opencores_0_avalon_slave_0_waitrequest        => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv,           --                                            .waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect         => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect,    --                                            .chipselect
			intel_niosv_g_0_dm_agent_address                  => mm_interconnect_0_intel_niosv_g_0_dm_agent_address,             --                    intel_niosv_g_0_dm_agent.address
			intel_niosv_g_0_dm_agent_write                    => mm_interconnect_0_intel_niosv_g_0_dm_agent_write,               --                                            .write
			intel_niosv_g_0_dm_agent_read                     => mm_interconnect_0_intel_niosv_g_0_dm_agent_read,                --                                            .read
			intel_niosv_g_0_dm_agent_readdata                 => mm_interconnect_0_intel_niosv_g_0_dm_agent_readdata,            --                                            .readdata
			intel_niosv_g_0_dm_agent_writedata                => mm_interconnect_0_intel_niosv_g_0_dm_agent_writedata,           --                                            .writedata
			intel_niosv_g_0_dm_agent_readdatavalid            => mm_interconnect_0_intel_niosv_g_0_dm_agent_readdatavalid,       --                                            .readdatavalid
			intel_niosv_g_0_dm_agent_waitrequest              => mm_interconnect_0_intel_niosv_g_0_dm_agent_waitrequest,         --                                            .waitrequest
			intel_niosv_g_0_timer_sw_agent_address            => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_address,       --              intel_niosv_g_0_timer_sw_agent.address
			intel_niosv_g_0_timer_sw_agent_write              => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_write,         --                                            .write
			intel_niosv_g_0_timer_sw_agent_read               => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_read,          --                                            .read
			intel_niosv_g_0_timer_sw_agent_readdata           => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdata,      --                                            .readdata
			intel_niosv_g_0_timer_sw_agent_writedata          => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_writedata,     --                                            .writedata
			intel_niosv_g_0_timer_sw_agent_byteenable         => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_byteenable,    --                                            .byteenable
			intel_niosv_g_0_timer_sw_agent_readdatavalid      => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdatavalid, --                                            .readdatavalid
			intel_niosv_g_0_timer_sw_agent_waitrequest        => mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_waitrequest,   --                                            .waitrequest
			jtag_uart_0_avalon_jtag_slave_address             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,        --               jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,          --                                            .write
			jtag_uart_0_avalon_jtag_slave_read                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,           --                                            .read
			jtag_uart_0_avalon_jtag_slave_readdata            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,       --                                            .readdata
			jtag_uart_0_avalon_jtag_slave_writedata           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,      --                                            .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,    --                                            .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,     --                                            .chipselect
			led0_s1_address                                   => mm_interconnect_0_led0_s1_address,                              --                                     led0_s1.address
			led0_s1_write                                     => mm_interconnect_0_led0_s1_write,                                --                                            .write
			led0_s1_readdata                                  => mm_interconnect_0_led0_s1_readdata,                             --                                            .readdata
			led0_s1_writedata                                 => mm_interconnect_0_led0_s1_writedata,                            --                                            .writedata
			led0_s1_chipselect                                => mm_interconnect_0_led0_s1_chipselect,                           --                                            .chipselect
			mm_clock_crossing_bridge_0_s0_address             => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address,        --               mm_clock_crossing_bridge_0_s0.address
			mm_clock_crossing_bridge_0_s0_write               => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write,          --                                            .write
			mm_clock_crossing_bridge_0_s0_read                => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read,           --                                            .read
			mm_clock_crossing_bridge_0_s0_readdata            => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata,       --                                            .readdata
			mm_clock_crossing_bridge_0_s0_writedata           => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata,      --                                            .writedata
			mm_clock_crossing_bridge_0_s0_burstcount          => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount,     --                                            .burstcount
			mm_clock_crossing_bridge_0_s0_byteenable          => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable,     --                                            .byteenable
			mm_clock_crossing_bridge_0_s0_readdatavalid       => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid,  --                                            .readdatavalid
			mm_clock_crossing_bridge_0_s0_waitrequest         => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest,    --                                            .waitrequest
			mm_clock_crossing_bridge_0_s0_debugaccess         => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess,    --                                            .debugaccess
			ram_0_s1_address                                  => mm_interconnect_0_ram_0_s1_address,                             --                                    ram_0_s1.address
			ram_0_s1_write                                    => mm_interconnect_0_ram_0_s1_write,                               --                                            .write
			ram_0_s1_readdata                                 => mm_interconnect_0_ram_0_s1_readdata,                            --                                            .readdata
			ram_0_s1_writedata                                => mm_interconnect_0_ram_0_s1_writedata,                           --                                            .writedata
			ram_0_s1_byteenable                               => mm_interconnect_0_ram_0_s1_byteenable,                          --                                            .byteenable
			ram_0_s1_chipselect                               => mm_interconnect_0_ram_0_s1_chipselect,                          --                                            .chipselect
			ram_0_s1_clken                                    => mm_interconnect_0_ram_0_s1_clken,                               --                                            .clken
			rh_temp_drdy_s1_address                           => mm_interconnect_0_rh_temp_drdy_s1_address,                      --                             rh_temp_drdy_s1.address
			rh_temp_drdy_s1_write                             => mm_interconnect_0_rh_temp_drdy_s1_write,                        --                                            .write
			rh_temp_drdy_s1_readdata                          => mm_interconnect_0_rh_temp_drdy_s1_readdata,                     --                                            .readdata
			rh_temp_drdy_s1_writedata                         => mm_interconnect_0_rh_temp_drdy_s1_writedata,                    --                                            .writedata
			rh_temp_drdy_s1_chipselect                        => mm_interconnect_0_rh_temp_drdy_s1_chipselect,                   --                                            .chipselect
			sysid_qsys_0_control_slave_address                => mm_interconnect_0_sysid_qsys_0_control_slave_address,           --                  sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata               => mm_interconnect_0_sysid_qsys_0_control_slave_readdata           --                                            .readdata
		);

	mm_interconnect_2 : component NIOS_RFS2_mm_interconnect_2
		port map (
			clk_100_out_clk_clk                           => clk_100_in_clk_clk,                          --                         clk_100_out_clk.clk
			mm_bridge_0_reset_reset_bridge_in_reset_reset => reset_bridge_100_in_reset_reset_n_ports_inv, -- mm_bridge_0_reset_reset_bridge_in_reset.reset
			mm_bridge_0_m0_address                        => mm_bridge_0_m0_address,                      --                          mm_bridge_0_m0.address
			mm_bridge_0_m0_waitrequest                    => mm_bridge_0_m0_waitrequest,                  --                                        .waitrequest
			mm_bridge_0_m0_burstcount                     => mm_bridge_0_m0_burstcount,                   --                                        .burstcount
			mm_bridge_0_m0_byteenable                     => mm_bridge_0_m0_byteenable,                   --                                        .byteenable
			mm_bridge_0_m0_read                           => mm_bridge_0_m0_read,                         --                                        .read
			mm_bridge_0_m0_readdata                       => mm_bridge_0_m0_readdata,                     --                                        .readdata
			mm_bridge_0_m0_readdatavalid                  => mm_bridge_0_m0_readdatavalid,                --                                        .readdatavalid
			mm_bridge_0_m0_write                          => mm_bridge_0_m0_write,                        --                                        .write
			mm_bridge_0_m0_writedata                      => mm_bridge_0_m0_writedata,                    --                                        .writedata
			mm_bridge_0_m0_debugaccess                    => mm_bridge_0_m0_debugaccess,                  --                                        .debugaccess
			SDRAM_s1_address                              => mm_interconnect_2_sdram_s1_address,          --                                SDRAM_s1.address
			SDRAM_s1_write                                => mm_interconnect_2_sdram_s1_write,            --                                        .write
			SDRAM_s1_read                                 => mm_interconnect_2_sdram_s1_read,             --                                        .read
			SDRAM_s1_readdata                             => mm_interconnect_2_sdram_s1_readdata,         --                                        .readdata
			SDRAM_s1_writedata                            => mm_interconnect_2_sdram_s1_writedata,        --                                        .writedata
			SDRAM_s1_byteenable                           => mm_interconnect_2_sdram_s1_byteenable,       --                                        .byteenable
			SDRAM_s1_readdatavalid                        => mm_interconnect_2_sdram_s1_readdatavalid,    --                                        .readdatavalid
			SDRAM_s1_waitrequest                          => mm_interconnect_2_sdram_s1_waitrequest,      --                                        .waitrequest
			SDRAM_s1_chipselect                           => mm_interconnect_2_sdram_s1_chipselect        --                                        .chipselect
		);

	irq_mapper : component NIOS_RFS2_irq_mapper
		port map (
			clk           => clk_50_in_clk_clk,                   --       clk.clk
			reset         => rst_controller_reset_out_reset,      -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,            -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,            -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,            -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,            -- receiver3.irq
			sender_irq    => intel_niosv_g_0_platform_irq_rx_irq  --    sender.irq
		);

	rst_controller : component nios_rfs2_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_bridge_50_in_reset_reset_n_ports_inv, -- reset_in0.reset
			clk            => clk_50_in_clk_clk,                          --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,         --          .reset_req
			reset_req_in0  => '0',                                        -- (terminated)
			reset_in1      => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_001 : component nios_rfs2_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => intel_niosv_g_0_dbg_reset_out_reset,        -- reset_in0.reset
			reset_in1      => reset_bridge_50_in_reset_reset_n_ports_inv, -- reset_in1.reset
			clk            => clk_50_in_clk_clk,                          --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	reset_bridge_100_in_reset_reset_n_ports_inv <= not reset_bridge_100_in_reset_reset_n;

	reset_bridge_50_in_reset_reset_n_ports_inv <= not reset_bridge_50_in_reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv <= not i2c_opencores_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_led0_s1_write_ports_inv <= not mm_interconnect_0_led0_s1_write;

	mm_interconnect_0_bt0_s1_write_ports_inv <= not mm_interconnect_0_bt0_s1_write;

	mm_interconnect_0_rh_temp_drdy_s1_write_ports_inv <= not mm_interconnect_0_rh_temp_drdy_s1_write;

	mm_interconnect_2_sdram_s1_read_ports_inv <= not mm_interconnect_2_sdram_s1_read;

	mm_interconnect_2_sdram_s1_byteenable_ports_inv <= not mm_interconnect_2_sdram_s1_byteenable;

	mm_interconnect_2_sdram_s1_write_ports_inv <= not mm_interconnect_2_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of NIOS_RFS2
