��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"�I.ͯ��5��E�����W�uGUګ3��'a��o%�k�FW˩���-��~X9��[�Zz���	_�qE�̟2V?,+d����ͣ��\S?�Y7�ZH,F0�)�DȀ��&-��Sr��D��҄
-�{F�GJ�#��j+`j�̾��Ҧ�U���w���ڟ��O~��`�D'h�}�.������j r3[oPٮ���LG�γ%���&Ϡ��~(;T�t %�Z��?��0�9��M��M\�@��@�k�B�)�>�
���*8S�!3[`(���E+�5z_ ��퓮O~90ڈXCS���7��'+����(�zY�bOK#�K���V����q�Ջe�j��-�[���֫�жLmGqOLanR�Zt�i���Ǹ�E��p�)m�"h�ԏZ|���죰�)�F��<��^b��%ذLފ�5�f�Ό�CJZ�a�<�y���/#���ݒ�!G����?��G>���l,�ŗ��ؓb�
W��A�I^&��B�@�L��� mD��r
�o߿���e�9F��G�R���s!h�j�Am6*���˕�5�gt����lv��KtI�r��X"�����-�����%
�Y9�%-�����{�ȇ��Z�����Z�&�?!촊g�= �6f��b/��D����L1���*8�>�����0@�z����d�m�^L˴7�D ��~J"_ϒX q5���"Z0��E�Z��C����򧟘�9iwt,�~����9�Z�0/�O��݇�b1Xm�x�]�Q�[9���~\�z��m�P���P�ŋ���r�)����H?M���E�צ����ɾ�:�'���$�q��^8��`U?%�:��B)���Z���1�z�����J�S$�g�ꬅ�Rst��a�9�Q���f�����8Qp�J����z�K��-2���:!�	��I�Q�"k;l1�@���v�
��vT@�[4�ﲧ! �t� ����T��w<	v��1SْF�N�oVÒd�`5��_��M�ƣ��]�F,l����B�ݪ�m͝1���[���śB��bo�����z��(&�?gܳ���5��)E��g�ZZr�H��KR��ңt�9��J�h�#���BW�֣��P5���$1n�Z#�D��]I����I�W�%����3YDC�1y��&���T�N6<ڿ���_�0l�j��MX��w����H��>{��ڨez�"���y�`��!�ը�D+�b��d�Ԙ.��*�_�-r��j�**����U��I,�J�ma��e Rw�O���J�{!�;�D�!q��E�iF�N�[�92!��4!Oan�Yˈ�d�������9�!؝�0h��L3߁����,��YhP�[}�.X�@~k.�/�=��#���*�#>��q�Gt<IRB�҅��E5R~�|6)5zKH,�[�;��a��b*�$�y��ߞh�+�-�-(��O3
҉b)���B����κ�v[ �ٶ�9�7`�g�^��O�q��ލ���dP?=���8��9��������GϥeyC.?hm�2O#|���l��<�~���ߪ�%G���dϲ�pA��L��h���6���󡋔U�X�[�_����:@���R��	�<��W��%��Hh?X�v��,��:�A�rd#|f&��#�WШ��v5c�)�I��D�"��V�Ӈ)p�S]���q3�=��k��t|�Q�<����uja���"FB��mi�h�<�J���ڤs�p��Z��5&���[��6y��z;pg�	e����Cc�9M��l�N/�>fGI̡xԦ�el����"�P�V!���)�+k�=�`�q%�^���6��k��9�x$t�q� e-�gd:�&�1�澫%��~ʾ��%�d8�5t�ޚE\���0�{Z�a���d��{�q?�1q�G c��PkN��N�m�k��'$�He�s�y�b�1FL<$ԫx��yo��T\���<p)�G;���J}�L�����U5_!�Z�!��Xu���׈nn��f�� �~g���ϩk�噾Q�e�݁|��SLr��}P�����2;j�&	�0���z ��O�7U.Š�ud%��UIY�9g�Y�i�✦��;Q���B�f����B����J�?��ί�q�@|%�P@w�:���R�#��{E�S�۴����k�]Q����q��'��?��,�<@�b48V��{��N�,���F!�u:��qV2�7���,�E�6��6��	M;z7,(k?F1_,;�Ũ���]�%BJS�V��� �1�F���x`�$�m��25@/ם�^����{���^�@�B�`6�����*�Idd(hi����H3�ŋnCCĚ�lͤ3��T�å�O�­���'8���P̒�D���J����!�^�em'Kf5�E�2'�D�?ȩ9x���V���[��9>�o�}���c�P|�p#dMV�:�U*XNN���%�A����̇�H̯������J���t)��~�_zk�!�3�<Պ��kI<���^�r9a�p��xP�߷q#�����P>W�@\=�uy��:�CD��J���\�^�s����`��3����3u1�^�Uer�1��@Y1�����B��]����gj�^�F�?�,A��T�k$��H����<y}�xj����k{�Q^xcV`g��8��`i-����YbE�Y�˨8�%���z�ռ?_$�I-����I��+�Z2"���o�����=Oc����Rٶ%��N�4��� ��g��z��!P�	�~_���{7r�G�ux^oZ ���{� �e�AqN���>.�T�a�?T��x�Nꨝ�n�.\tXl(}���i֮F�!����_��)���奄,�&�Yׂ���	sa���L//�Xz�CMT�10?�:��C!i=���Ptv�ܓ�]&�H��>%�Yyr����WgC�l���>j����X���J�;Op٠*e�"��W�Mi1�ix�� ��������-�Գ�C�������g}�&��nzY�����C�>��6m)_o�x�����?Ϸ`�����:.�<�h��P��^rwoT�w�-L����k�Z�}��Uj�k}�4�������dc��4kwf�Z�r�~5��pXΨ��k��8�:���c�|����]^)�������oB"�-�.�40�u�ڑ������[JV�f �J&�ڄ��o�� ���2��y��JZ�m֗���x�z�`��˥���h>n:sl~+���8#�0|���`$*��$:�<�H�_���Q�E{���rFna|��Q�3��f��}�j��J��r���#AoOd}���Hg�X��CXa�G���x��~��?+]��߂����|�d�H���]GҔ9�]]�������S#A̕7�t5)���s�t\�-��a�n��PL��1;��cw�9#̄���Ww��HP�ϖfCr�) �P�v=q�o�W�@����DN���
H�XSD���Ǚ��L"~0W��nB%�G���Vߠ�#���?F�N�g�K�ߗ]?η�Ai�m6�n�?e���	��_-I���!p~�'��us�N���L3��P�Cыـ�������&�"J�Tާk�kHV�Q�?�{?=#��Y"�.P�]��t.������De�카��	�e�e�j�gٴ�e�s�2��Rj#Ρ��"��av˝ë;N�7+m�O�!��NL{)B��F5�c�5d
Ӎpf��Y�U p^Yp���-���b0z�n2,d/´׽jB~���,��|8k]
d�@2<x�Ah�f�Y��F�{N�'�����-Q*�y"+���ȴKӨ�A��	<
���E ��Y���.ק�.	���� c��8ّ	�G.��S?)p)����B2'	�OM�@tl%13��΄�eq�8���&7wn�4ξ"��_��)P����}0��H�B'�t����n���}"��zo���@�*t��gY:ܳ{f�0q=�-���L��5D�En�?;�h� bu&�-FFx%����\�9�
�^��i,<�z�q��np������?���o�߮~��CpJGC�j�+Z�#p2�1����N��J<6[�X� ��ӡ�������6�D ~	\�����f�r��,����	y�i���j����f�������}���o�4��@.8A	I'\�q��ٸ(�������o���#3�A
�1�Gq�U�9#��	�����`������G}�����H:0��pM���p�����F�����u��O�d�>9�F�-<�	1�6�
#�K�b�Z!�mj�04�yݖD}�:z�'����\0c9����qV<�H诎��x��&������g#*D*j(�cqoڰ����F�ۋC� �����R����OKB4gUU"ة*��	���D�N�ҹ
���ᔉ��#�ֻ�����{+�\!h�i�[SQ#�w�Ѫ�Y]M���6�y���^t�Kw���%y��)�"�j�Ed®���B��7�<�.�@��
u� �Q�Tӧs�~��, �%�F�A��#�*P�ϧ�f���ɏ�yҾd���(�H|�$�h��PnQ�ܸ^2t,��L$�f��ja�$-��k2���]����~^�V8�WWN�t�*��B����a��J�S��,2*��u	­� M#I5M��^���w����͋�{�M*��_�p56A�І�x;��9���.���
�.��M��>�9���=��{y�OY�-^����/���=E��D��8�h
���u��.sV�@��&c�.DM�i�j0c�B�w���X�g�8F������ffwC�R#��,y��1���-Pc�W�����i����9���*Q��3�n_�;��N�hty��2��c���L^�
yg̭�-X�:�Bz'L%�{d]�����[�l�F<���!�j�����__t'Ⱦ�m��{��8�.�B��./�>���T��IԆ�o3yQ�`{ҋ�|��׆��m"s3�7bǓ`�t9��K��`�KZ)K K�a�u`\Ź"����2?Їt�]�F�5k��hS-*rar<#�ݷ��{�*�������E;�w�a_2���ۗ��ѳ!�+uA�-�@�+\pI �rW_]�U�qUA�fgՑ���1��ԥv�UјMK�/}��T;���e��k�]&�o2���=!�s#�_,��|�i`��ᥢ2��@�b89��q(
�%��ӕ��
��1�6#�5��V�E��!�5[��W�����ʺ����P���kS"�1���k��N���li^ͪ�����>��t�s�!g���Z�M�B�ɻ��Ȕѫ�J#�KeL�^��G��33�˚����gK��M��h?��q�Y"̞�-v4�X�ݣ��&