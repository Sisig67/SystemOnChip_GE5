��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%��}:SJG.�O�� ����ƊBZ���=�Բjr�E��d&�녛0���vS� $X��R9%�zt���\Vf	����Ķ�����]���\b�ܪ�F˚m�K0�h�:�ȕ�������n#~l�0���<WCYХR+p��4��@ѫ4Oa����T����K�T�ā�Z�L��� ��0�y���j�PdQCc`��ϋ�ʤVD�\�� �8i��� �z�9����tPG=����Bڽm\6��f��]���&ԥ��n k�>OY��V�ԧ0 ���Ӛ����xb���Sտ�RJ@JγRN;�Ȭ�n2;��x��+�M�<�;�2:p
����\��vB���#hJF�S�]�}�D�C�~E�-BCH,�35:��l�
�b5�.���L��(�#$�+lN\�ǔ/�*4$l-��l���!����L�Qu�q��n�W�l����t3wq� :��aYA�0M��%Ҝ��;��6oJ[T�^�q-��3Z��=m��r0��?����4I�>k��=㥲��uwC��>�.���~2_z�4l��}��|��;���z�Ž@!��/��������:�FǙ�_�\n|�D��\ޠ�)������IT�Ƚ`����r�!���g�ĳ�	���TS_F��v$Wp��v0��)������W�7TBr�5����j��+����<���ʤ,&P����`k�U7���ΐ�G�<K�э�>��@!:�v2e@T�DR�$Ci�%�O�-�HvX���eUns���	X��!�3����Kc�X���ͅ������E��z��UV��nx��nX Ư<h5I�ǚ��BK��͒kƎ����4���,�,���~�@�j|UӲnU����yAn�L�����t�x���ʡg8@�O�hL� "L������U�4������ohB�c��rf��\V`�2�����e
���eBI�+��߅(�Lsm�F2\
�磪��!���Q�=���{$c�����N�0�g)	�m�c���اH�0�����H�� �n����]��,��欇�ωAS�NT^�|$��+��Н����(Ϊ�������n�1>�C2U��ՑsX��)Y�k�Q>�˂�����a똊t�]�[Zq�
e�;4�Q{������g˙���S�+�a��މ�o��DZ�S!5�Y�"I��x6&R�Q4rE=`�b~p˵���tj4"���5���L1�}\��\�)y!p]�t�N� ����d|�k�ʨK�7[*Do
eʽ���V�������k�}ԟ��qX.�
l؃N��_�☩N��<�]v8�3�(��	LGQ����K:����*�{���t�2�v�F��8�i.��c���ʗB= !��d�n�seɉ����kb�M�#�ѹ���>�y`��r�Sσ�h�m��S�z���}1�` ��ܸ,QRq� l�pq��/l-.��V�Y�����"6�����k����\�=L�:qo�w����&C�>>7a}�!�����6�AG�"Ju�Kwٽ�%��U�mCUt%��=�m=�Uda@30Ϸ�)?_��l(���e�ǡ`\x�C�Ug�P�e=�|�z�����x���&µ{�6��镥xk��Idoo�˳9ca�*1OM.��8�o�e5�K�Eo���MѪ���j�o�̪�ۍBK�Z����_f�O���@����)����|+��d]`
��gt��N��J��p���y�-����TQ�D[.M��,����fݣ\l�ul�!�T��"/L	"1�Vh�1�|�q���C���y�K�֧+�^��T0�l8m�/$P	|$�249^ꜷmcm���<W���������~���:�{ ΧPDFc�[����6���$˥t�D*��NH�7�v��j���+�G�f�d�����hL�"�Ke�FM�R�Z,�c	3D!��/�]�A�{��%I���k5�Q+ー�q�i�������sA͚U����?�oBo�� ��9z��V%͒x���>ć��bp��^	535\,���2FdqF�o٣�=`�����d�����	W��Y����K��q]�7�%�o{S�� ��pa=�����ƕK�c(����bp�|�"\�ڴռp���r	��#��v�q���� �ޞ#��St�'bY� 
��\B��v%c���r����(Q���5p�4��5�3�S�v�]�Jgi ��80�:�tM^����\�zXt�ϑ�qT|Oe\�	E�]�:٪[�o�~�nmca��r��c�M��ڰ�+� ��ɴ��|���C{�&��m����T�JCg��>�9i�U��W�,_?����%K�C����P�����Q2ޘE���M �����2�-���ח?��\�v;*��Jt3�p�8U+���|W���1��7��A�#:I�=��P�g��*A�|�JjB� kb�Ӌ;!�M��QZx�E���<:�C�+���:�?���`,
��[mMJ�Z�����ڙ��̓K ���QL�v����i������)f`�a^5^	�\���'�y�F�U�pCb�U���QMƸ��u+��-"S	m�G��D�wb؁�e�������@z��6!P:�Z�-�6���&��M����U|ql@���Z�ۇ��ݭ� �O��c��]8��Q@悘��oe���4��[2\��M�Q'ݵ�3S�Us�'>�cN������3D�8h��tn��?T졹c�i���u�ڀb�&	���)[�n�uZf`����x���ꃮQ��`-OUj�iS�F{V�wg%�����ߵj"z^��M1������-���"_n�^s� 6"sH���v<2�C�"���������ӊS�d�Z�x}S�u9=�Z�腓�L�����6��~��Y��6?���n�2��=}$d�W�sx��
�@��%����eHש�!�ݐ�+��#�Y�nJV?�<q���dD����	$��p/qc+`u:�+�#V]�@�t}9��fQ�� �$�-�j�G�o���a�C�K���(���[M؆u�=�m�΅q����\����g<�1hmy�	B5$��>���7}�+����U�4Uz�>..����>�k��F�h8��{��
����S���d��i�i�`fR�<�[�w�*"*G8�4q�d}�Q]���x �a\B��C��;����!����=��$L�j�&Xet�f:li�
��QF�Ve 0a����zYPt_C4������K�=�-�X��ڤK�[�5u<D|ȏ\�ȩ܍%��W���� E�eI��N�U)���·��y0����+c9����\��Sj\��i*w�A��s%2/�' ����d��*N����#$����Aޭ���>�y��
�N��0f�+�zy����:���U<��]U�vc�ގ�V����?Bsi�z�ED���,c�/��9^D�/���D+���M��n)�������&+�則tt�!��������v��L���	�('	\�#�-wS��2����X�p��Q�������uK�KkZ�
\y��{�1������	!(�������M�>�+���WaX�z�	};<�B��O�1�gc%z�ߩ�b�ѷN�����4�^Q�f��9��O�HP�\�x�!��I��T�PM�x؏Y �(!��H`]�-�/���]`��36����+0��r�h�%
J������|��y��t�"��lg&�y���0M�v�镓�S�g�%KԊ�7�T�X���j�t��������4irweb1����	o"�*TJ��}rS�/p�����t^Z�!��A8!��@��-^rP��u0�N���˧DZ��J'�v����֞�)wԘ��.����'01x%N�B�:���Ga{{�ɐ�!J�(Q��_L�s5���u���kR�ҝ_�fF���C&�aN�(����3��(=���_��ȟ�-��\���=��ǔ���`�.u����Ė�R�.����\�t^>,�V��=�7ke2��Ipn���t�]_�6F]���D4�As����
9��bq�D�'�Z�/��O�z�TR���Éy����R
i�3vz����4��rI�s7[��E�%:W�F�h3TЧ�J�HFIt����J$�V�>.�O���̋CG�k��"��N�L&��e��26�ok����&��e������x�Oދ���>�6N�k�_ٽ����O<�}��,
w�_��0�ђxc��Ƙ�]z
V��6�c����.fP\�f��I}y(��Y:/���%���@�6�U����V��!�nx��&¡���ͯS`�q�>
#g�8)��y�˹x��S
܍�<����d��T�X� �w�l�ed���zW��Y�\d����݃���L97?�3�H�]I����+\ź��'iV?����2\}��)�b"�9k֞�C�Խ�� euX��6>����O�"�%�v�	�L��\/J�1�*���D=��A�VתC2�1���f㳱� N�Q�(�t��0Ʉ@�u�5�K�rd&AH�
6y��[��f�UVrY0	9�W�`��(Mv�K�'������ɶ�72Õ2�6���)"����Ґ��ܾdݻ�;�cI��n�7�B�fv��I֭���߫EĦ��cദG:l�u�͠��Uz��4u���~����Cc4��^�2J� e=�H#�օ��!�K����?=�_2R�l8�
%�<����R>^��n
;���T%��}�G�o"���U<�mۑR����e�YDn>w�\*n��X�wE镣�����k����:��9*��&N`k��SP���� -��0>=�;J��3�,���5)J�H�B��z���0'�Q��]��;$�vC�Uq5�w�U/7#!�2L\fݾ�,k��ʬ�ɏ��/�Q�*U�`J�{i��
�kڵ��.(p4�G�n��C8
�C����'��B��,�s��ܤ��F� 32L��٪9yŔ�����r}�>��Y�z�Z�ֈ%ڞ���D'�etw|K�!W*CTmWG�CI��K���i8�%�]�䦦�մ��q2�ԓ��ƶJVS;�qT��������
�{���Թ�w:�R����9 �P۰�v������2!au��X�%8���c��޲l7�)-c�mc�m�[�^<?}�M�z�f�Q�s��25N��+�h�w�\�FQ46<�:���\O袄Ńwm��n�fM��C�����>�K�}1Y�>�ZאY3�U/C�奈b/��Ί[<�VOf�s)]�@�=hZ��v��ӳ6��t��8ҋ�MH��Z5�R��*�j��O� �/!�K=�d�ްB��eZG�Y�i�A,��M�W7P#���$z�}�N<[�$�?6���D*�ql=$�\�\�M�mj	�����c��&w�yZ�:��E��D��5K� �oU�H-ީI���zN2�!���ӐUA�?�:��$KR����.�9W�����j�$P��"Yf�}Y��)�"(�2�<��[L^'��+
��Ϩl�J�[�ǿ�"R�<�8ϡ����.ļ:Z��B��:k���S��eQ�Q6]%�
���l����Ͽ&�L#VgL.��M>���Jy@�&���|����(�^���C��V�2q�E����X���R�3u|!,��S!�w
=!�?T�{l�R�ME�R���,�l� #��gEʏߣr{��M7x�'�R�}(�V�;�5�y�0���Y�����!�n3;1��;UT��Uv�o�&����W� ��͋�#��,����1:Ǭ��	�Jp��e��//.JE�����;�w�|���?61�fa��d��5�BEw+"s�:{��ۻ��㞑͈&���"�6ҍ�6�*�*�샼c�=8�(��xd�j�g3�h��lű�h���oO4�+S?{|9D5����w��+�V��5���a�k��f
���5RZ�!I��A=��ck���Tgg�USӁ�x5�q���l�	I�"���*��$&�g}�K���B�y@䌲�A�	�S�A�I{��/vȵ��h43W��Ċ�ʨ`�%b�z����GI�`�7��H�<��gA����H�d�8�}I!��o-�ק����b�,����L\]-�5�z4Y2s����������.�l!й�������"���W:0�=�Y���ik:��F�~�#@'�o�~&��'I���1�l�Š�<c�0�7�n�b�3�9C`�RGD�p
��?���[=����n-)�j�q+��Wb������3� �Tm�~3,����^�g:X�zp�E� ���	�J�iQ��wx���l\bC!�u��7��&`��.( �~�c^�f�!��(�� �
a��H4��8b��w�\}F�w4�`ؕ j��� ��l�!����-� �1�$皦ս�>���	͘��a�j8Ǜ�*o������mq++)!���t,3@/	l�e�!�Na����)&����S�N\�s
=|a<{E���9)���o��� S��6������)���-����`u! ��S��r;q�"��.�q���B�Jt��r]���ws�i��0�ч3��唳q1�u,����ڢ���Q���U�^�Ln	,
e��e����	@��Ha���4H���?�f���v��<����a]{g��d>��g����LuC��xv���1�U����l$��%�v�@��,�oP��t*���<f���^Nm�d��3�$P�TbDq�!��L��n�-�*��0�v��\�W�m�bE��9tvvHu��d��Mpʓ�����?�ڶ���lQa���é���8��^����"Ҥ�j5B����X�Y�֪�<X�ˢ����Ju�yho��n<���iV�z��t)���W?�'�o�s춏����i_6:�.T�g��~��OJl�-���G)؝��
�n��a1J�x��6�C�8�TZ�N�ȣZ��i9U�p�o�(8�����;.S���|��\����g�������4���3'�Kb��A�}�B�VU�:���)�Zi
?�;>1��sƞ�ᲀ�녆?vxC)Ęl���0���^Qw|U,&֜�2��dt�Q�X�ʐ���ݣ�n[PQ���LK��l�$-+sC̟�W�Z����1v6��Co��w's��{zz�����tx�g��d�M�Յ�<٭PN"�6٘�A��tgyP���x��q�&('a��+�; �$fG���.Q����9�����j�g|���;�	"f�[1�T�/��q���#A�^��sAI*TG����A��U/�|�4�5R�+�>�0��N�mp�i�&罆�ݜ[����T��5�����0.Z�M�k����:A_��zzѩb�?��NS�f���o�������>�������E&�+Yr�Ɩb#|{�kS�VL�L�� �R��C=����^m�x��PE��~�0�\*�0�꺩^�tx͐VAe�Z��m0������W���d��msqi�̺1d���m�Z4�#��
)���ߚo��Zx����Y .�~,9:�];n�Le�ӑ_=�6��#pi[V�h�O=f\`��v��h��k���m����-�h���9˷kN�dS'w��� 2���g���KS�)��L�t�G�-j;�D�؄"���3�_�%v%u�Z��Z�{np�}@��E�*�sx��p'�'�6ɂ��S�����쐆���a�Ϡ$v%H���Zv��*�(T�V`�洽�z�Y�wm���di���m��ǔnf�<η-�����8��K#��c�G��R��u
?�z����q���R�iui���y]�xۮ?�O?�8�R�l�v�ëYf5V�Ű?f��������P�O�I���QP�Z�ȏ"^ɋ\زԖ�$�Y��3JV�ٻ�x&�(��w_#$ehoI@����~J�QY��ї^�Z}oXم�HJ���ŧ�2� ͐�n%J<�PD�/Av��F�YI�-�((��Br\ �� �ޝS&��) ��P�쁳Q��n`�)VW���Z�Q��V�#����1B@��f��\S�;-(��lq�y��p�-O�!$\(�q]�~{���3P�8 n���3 ��1)�6��U�Ӵ�F����G̭C��?B�abTe��r+��(�]B�nVs?�O�X�3�󘔢B.���"GܙΔ�$wr^���1�1�)9�W8�<D�O�YnŃ��7��n��L�]|�>I�q��m�VcMן��,��6�v[��2�kܖ�=�<$�"�H n�?� �G=� r��{����	�z2"�1>��/�zq~Ӏ��58�J�@u�%�U���i�o�+o��2�'k7��aK�	�)����)��Sp=��Ѥ�APB�5}t�~� V`p��:4�l �6^�;�_��	��Tǐ�I��'�/���p��5�Ě*��(8�2r��x��S��%PEE�1X�r����\����<�ӌO@���Ճ)�W0~�tE��0?������S�z��4���Π��,O�6W1m�GΆ9-�OM�Ny��	b�S�`���7��1q��5�7fB���s�8��A�.۵Gs=����̗�N��5*����YY��^���5���?�� 5P;X��5���:G����Ka-�r�%��4$�v~��jA���5!��l-��Or�$��b���?��'���k������_����E�$:Ը�ZH'�i!}x##��#�/��(qbT�%<�?d��c�3������X�`��Nj	�[c�?�>�Ώ񥋙�L\'9B�aDywX��Z!0{H)�]�a�(�p�'Gf{,�C���P���u����l��/��YgC_ME��@h�(!�{�su��O1���ȁ[p'|Ԣ��S�ג�9���>A#��H:N/���Esf�&D ��;W�����dd oe[��j��^Qޜ�X栩��Z�<I5��b����c�%�(���_{X��\�+����U��WL8���~����<�Ɏ��AWA��q�Z���zꮩ/@G&f4��wX�I��8�����k�G��:��%�- �v�,,�(y>�B�j,�i��Q,�\H�2��|���} ��:��b���YH��P���N��Ԃu�Ar���cw��*�P?]nD�'8����.�f�u�$�B�K�	{�l����|#�H<��I�)�ĳ�3�>�v��Z�Q#��*�TIM!��D/����?t-�s�}ٜ��[ge�v��� ��+n�2�M``��
Hi���(~aZ�@�gP*KQ&u;�Pn�;��0E7������'��
���ܿ���ُ���d���9.�,�\V�"��gu5.��~l1;Dt�}��:H֣�(V���u�nk$l�a���2st��GhY<h�ü�JDZ���(%N���eX�z��@���.A[����^n2]<�5��I�j]���V�;f�'F6VG���/N�HY��4��e�~S|â�RI�H,�$%���<K|(�0�VÍ#���=Ӝ�
�O��P���_��z]ε����������+�\�%kVq��e(Q�wZ�0�L.XƠ|>N��:%�?t�^��]'ۣ�S-GЈHp�\#P.�!F{�a H,{��p:�x����c����]YSwd���g�o���2N��P�:����lS{.\�y�}�������&��+���e��h)G9s�#a;����P��S���-u�������8\�����������M4������((jr�YKW��W���l4��ZF����wP^V�I11*\�W������}G�ʼ�L\��8>��G�ҦS������'�M�2Xݽ	$�]�Z�M�+���y�D��(�� �c�b;�D��e��VP*�S~L�����#������#�?V��=�\4���`�>0�0���½�t[� 1�Qa�J�e֭��o�,�Vtב�/wLC@��j���y����pe�4������6���9����T复��  $U��U	!�%lI�˥��֬�!��.p&�>>B���z:��K�l�YO�Q�U���)S��&�u;n�k������4cO��0��z\�/eϋ*���Pj_�1g�*���p�Ψ���cId��Y�����vh������#l���W%k��5��{����1�ڶ�5���	>g�O-��$T�N����6�U{��l'�u���L���*�u`j�-��/�2��-s��2w�{.0ړ��L�ĲP�=N�Oy�K*��<�'ڹ������=��p4V_R̒��.��ٵ��4��+�zNۙ����z'�2�j����R�]�@�evgAڿ�V���h1E��%7���5����-A[�f#����~��b!���R($�hn��#�S�w�Ds ^$��� e|W0�
�8���>��0�9��I��v����X%S�����ްBnI0;�	�8��	:11�c� �TgJ~�/�%7�!zos)HW�A|OG�^�Tmܤ�bk���VF�#�	\�Ҧj弗ߤ�p��$"$Y$�½t�`���2-��������Rp���*�2E�J���&�t�@8���'�_>L&�c����M�� 4�F��o%�$g�S�W�Gl�&�ϝZT�+�?l�����!��_R�_i$J-1@D�$�7M|��?���2H+R�"A��q��kG�0�u�̣|B��v/�r'i>5mL%�C��G�5���@�SfȕdjT��_�����9g=��Ŧ�V_g��7��&V����^�0Bba|����Mq��WZ�;�f��N���k*����b� ����'D
�DĦ�O�<<��$��j<	�r�����Cr��拽1�v�TW���ys;���lG헙�0���$ S?׵����Na1�D패$D,���_�P���ؒsR����,�י�o��`}��yٴ��N��0��/�3������8���DQ��]P�S@�Ĥ�F	[;�:F_t�"�A�P<.�|Ĭ�!�o6v(��l��J�Mg�۩t~��^��`}��8+�+���JK���~�۾yS�K^)�O��r��q�13s�,nec�&�.;lI���k�AQj�'�Hq����m��Mό��K���(�K��'Y��2����\m�C�z~�����8�Կ�¬��x�Uߡ���CB9�O�����b�����3�4�h9�0���?�0�||?.j��S^� S�T�P/Ѵ�r����Eh�=��䐺"���كj�������Ŕ�#��(\_�Sv>
�M�HH�V�.�����I����W��\6LCM�ug]Xx�q�jX!�Z�2!CN��t$e����� ��Z��?�����T�i� xqW���#�lS����e�h͕Y�D�"��R���r�n��-�A/ ���֡�&\s�(�4��yB�z�������������[�?af@i�C��z)��<ʱ@���Ф�pw.~��_��+!����
Kӄ��2�L�way��/���'٥�"���80s�dg���Qc��/$[lc��<�&M[x��LW��b�a���^��/�wb:�"�����+.<���1�3���Rs��hW��ccD��.���>��G�;R��G��<V�PGp7�P��%��Jw�ͦf�M�b�/�w�{���<ƚ�HSٷ��r`I�"����������*�%��n��T,C����mW4lv7�w��P�'/_6x�[�l��a�$۬�6vIu������Ku���V�o���k?�!�,p�!�.mP�@z���W��ե�X&;r����~���$����.������R�XB���>O��9����(�:�Fj��u��+f �A�0�-q�X��v����_�ki��7ܾ]�-��qX�
�q[�/��i��$ם� v�z�Me�#�m[��<2�kcޗNTqy�N��\��lG1!�Pz�Wd�ʠ'1���
~�F\�jG��Z��~ބߗ��T"hxD3ܟ����ד�u��ZJ���.�~�p����P��ô�4��4����(Ʋ���H�6���$����z�Aad�L�N��Z�s��U�4-z?��q�n�O�*�Uʥ{�!����2��@
�����S�y[y����-��
�8&!ڨ�]���*�m[��4y��-� ��n7����FҬ��_4�w���r���s���],y�n� 3B�os&�����F; ��$,�|�i��ZD�g ���/\�ӷ9��������0�qOJp{:�[���
�i9`��H���}��y@��h}����������ꩪ�~�@B��a�qO���7���ibQn�}aNFTp.b�Ҁ0;�����)pԪ������#(�����@�e��6 ��
Ҝe	rH2���$MKҫ�$gj�3+�
��|B���uk�ǶQ�^&����S���-X8�.^�-}"9 �d\��U,Lb9��vc9swڟj1 ��^���A�@�m�z�i��Qp��tB܈�R��D�P0j������T����?ȅ��j퀉��h9��~ �f��Bɠr���Xz����=Q�������%��Xlsd�@rxHI��b�C�\�}���*��@б�^��1O�a��4�]�)���l_,K�	�JʝK��"<�$�a7ŀuk����zdc��[��8E�2�gjBtȦ%���B�6��2����K�[3잾�1�G,M�q#:���̆k�Sá�o�jN��y`f���N� ��Jf��U�wZ'�*^��%"�D����:�Aמ�X���i�4��L�	<�?PX e2��x�oa�JȃL��x��bs��Z��D�I������<�
:r�4S����݂�d�����ȣ�;��W S0�dʱ�V�<t���ֱI�H��,�m^�b�{! Έ ��+Bώ�_�	&q�j��rzbڪ�����de��8Iwp��>j�a��T;�+�|�Z����pw
�<��L=���0NRk���g������88�pk��F�j?5��1ڐ���fk�����`6�eM m����G1��;�H���I�E��ooy�����K�Gֺ�ϒ������O����F��%��
ʼU��z�S'��Әs��@i�A�!�vm(a��;F��#+�r��©@��7+{��kWFH�4H*�*r��p�.]1d�]PI��X.	�&��lo�2d�f��E�'Aker����h��,|���1���+�ک|{��_"�7�+;75�eIcj�m>�s�'��zw����
�A�7PY�nׁ�FTa�'[��AY/�@��\%���R�-'�ȉ��>v?d���V�*f�b(>����v54�^��Xc��7����e����v��B<4�3��0��Ē�7T/�D#����:�m|#�<FG�5�8��sY�� vʯ��r�P6ߐ9����|G+Ll��B��ⴅ�Ek�K_A_`	��E�R�?"�b�4�Ͼ�n�#�V�Q�@8�Pt�F�J�]���U�>s�h���fz�����֏�@�e���67-BW�}�I
D��N���-�s�=�!u $�tq=g^�F?SJ>���?`��[.k�CJ0{�A�0F�� ʘ&O,��8y�o��h>��ݸ'�ǔNDM`ċm#�+��W���5x�H�8r-s��5�;}�pQ����_ȯ�U�2����P=� �/�OV�4���îT���w���̆�P.���)�k�	�nO�N�<�"U������+Tb�/"{Ď��^5fj�aՈ�LDkP��J�@#�ՙ��[_��:+�	&��p�j}%�|�2�	�о�+�����_�ûm�i7��"�4����-��d�����W�C���S@(�f@�ͽ�I� G�*6^�2�.0ӧ���t�pF=#��E`K���oD���C�'c�8*�XD�'�����Fk\Qr|P����ޟ���9A��F'ˏ�[H��z*r��S"��(i ���}5��(_G�<ΔA���#��9��S�UI-�:1js� ���V��3U�ܨ�C����qd fN��m�e�h!awMt�&Rw����o�w�l�f�����3;nX��P)<��W�����8춽�]y�2X_ ��_��.�5�9� h��#=�/8����oy��uY� �d���2������0��賈�]T
�hH�j�2lxЂa��ㆈ�:��.�Y����fS�J��0K�z9~�NX����c�pߝ�Ɓ�9�.����:9 =�E�-O�[�ɼGq�/"�g\ �`sO�� y��	�y�DҔ�:��%˰9mc6װ?[��$g>��;�{�~���5M���K�]I�Kŵ�0;:�zFZ	5���3�ԏ�6�y�>m��5�]7����"�&�Q���ΰ瘟w{&
��Ewz�ܲg�ф���H�55�/a��|���D'�]��<���Q�*��L3B���Ey\Z����	�c6ȭ�,�N�#@$»����m���C����z�Z.J�<�����0x)���4�k�I�j�[x�`�tp ���9D�f:z�x#��X�(.�'�SB���6��(�P�pI��a�(1镘��k;%ּ)��� T~>���F5��.͵br[�����˓�YA��H����]�X���:��Q%��~ �C�)Q�j��: �L���7�s�[K����Q��k'�a�+�7w�kx�:v��$r����}�#�@�����¾��om#f�]��[�C��KG�j��^��1.߇5�q��F��d3�9 �o�Wf:$��>�(1=���J���q��M�6�?�����������S#������CR����D� ?!���v��L�d�
-��pܺԌ�!�����h%�� 0�����xqr�6|�����A鐑���D|�V�q�������.�%����i�'�Ĝ�dj����,$��M�+"���P�!����5�H�s�/%b���1�z{�}6c���} ��B�a�!b�!����s:O� �t�8�R,�0H�>1�B�FEα�t�|�̢+���M��Ș����Lt��K�ɀ�KX����sB�_����!m ��p�d7)�z�� �Õƴ���\��ޅ��t�қ����>$�GhXJ��ذ'����^�f�3�'4�Kd�1Tfj~������TǑ� �,�2x��yH"W'�B2�)�+����c��>��@�-S����[gO����&Ι-n��+P<R�-5�C�>��iW>�4lxzU	���N�3�ëφ1 j`/��/��;V��*�&��������"�<	��^*G�|,}�� ��gQ*CR��#�k��;q(g�iF�;CC�ꥫ�M���xe2��hq�s�O8rg��$k����є��в�̨]	Љ��఍���J���f�*?���7֖�p��#���`�R��D�^d��`�m'{���G���I�\���������7��2�s�ᰢ�L K�p�0a7[�e
����|�~m>;� ��K�h�& �\�����x�=W��I��H�y�p�4!����Ē�\=���F�:�z� ���ʻ���h�)~�/q������N3���sfq&��́�1M�����G����|J!�/9Η#C�kq������4.3���"ײ�/	²󟭚�/QU�=--�O��
>ƿ�əg0c{�;�����-JϿ�+������ӭ���ϰ> �D�g� �c[�=W��}m��qS��a@�0��X�EQ�2��Φ��6��:4iBT}K� ������?B�h��*��|h�%��n��4ӿ�}��笟U�U	�q��1��u��J�@�R�q)��Ƥ.F/���AՑۚ+K��Ha��\O�W&���4�Aݦe�<�Ξ�fBaI;�5���&.�*��_�'�!��F�|J�f��'�i�(Nz�^�Ys�Q��T��E��r0-g��ox�}�S�c��Y�F� X��m?Ls�̞�z;��Vi�2�������ކ�7+c �uQfd,��V��f�c�fc8�{,򌿥�ݺ ��5��:}�K���tc[�%�QOU�]�J!Pc�M[O�+O!�3��x�N�J�|TW��~y*b!6:�>L-�|�B��T�)�0��k.�I��՗�q !�A4�C��^�n��O+-����θ=6Φ���_{�/�0�I&p�ݙ�%{�"a�k7rՇ����A�F̵ٚs�L&�2��I�n�N* A�ώW�R�i�ȴE��MQ �}f�����3	Z��^J,[�;�wp�ݨ��9�&M
��o3���\��[X���}���i���+�m�cL0n���Ta����;
z�5$%���,����{+��]t�Ln8��~֩+����$�9�X$�>�CG581W$<<+U.��v(aढ़��;K�%t�@�.��XL_�l�B:ZGW�E'w�b�r-L��'�Qe����i��]� ��yl�� t�%�-û�j�����s�anh	q�35�F&�<,���,ԑjI직P �y�-��p&�	��� �ө��ς��6z��i�~��/�Ɯ�Q=[70��.h���z�? �D�Xʓ���Fn x�ɿ�[NE�)�2[��7�~���� #��W�	�j1��^�9h��+J	<[!y����D���d&�Ԋy�2�����$"V��0l����(��S&X��-�fd���
]��c�%�xc�R�a�!_��'�1�1O�lR�~�_p�<��N,�-�]��q%�l��i��-�|Ch�r(ۃQ���BP���g�nj��`�~�ʟ��*���OΝ6����YjR������kG�wb�P+���g�$(��@�Ħ� �ޒ`��^��X8��̟lk_���>�wO%/
�a]��Vބ�?|-`�G�y0�f�9������+�B���L��%@L����Ե���v�>G�*�Bf,y���x؂��?	�2je��y{�ވ�@a@_%އy)�:Np��502A�jZY����靉"z逸�Ğ0�����_�9]���|:�F������#�c��s)k�$X�	Ե'�}�b�{��kS����������$��ư�f�}����f1��4���f8;����$z��0"w�����JP���h ��'x����_냰)�t��O|�	Pcde'�
i�d�k�Y;ߡ�s���R�-������}��y�[FW׿~��9���sb{���[ʒP�I,�%>��z?� ��-7��*��ۡg`���M����������9l�l�$���q����N��ۘ}<�A�&4s5jcB�� �Q��Fҭ����n)b���p�̬��Z���ڡ��F�yd�D��w�g����X3/�̡˕x��ubF]���2_9�4�aq��㑕������E����W� y%0��,rM]m�Z�yK����R���Q����tP\)t�P�_�xܛC�Kyܛ��Ko�y1�FO���}�yƱ��|��B�4��o�j�q�s4k�(�^��Ё�/	̿ŵu@J�(`,@�X��فkZ��+�k�1^�¼���ý��XV�("1"J^2G|�"����[��a)�`F�;U��Z��A�����ɞCۤk�~��8wzc'�#K�804���-�M=HZ�O�`8h��(��B?ȞØ��0# �t��pS)B�E[g�:���~�vx�B�r��[�/��Q�<Z����$����4[��\����G$5����=Rk���!G�X�
��i^�@�-�sA�$UM�\:ĕV~�)z��3EI���������UAX����V���J�lpgh!�:�����u�|Y��\e���MQt�7E���L�������zֈ��5f�ΓF�"6�������ehL��G�?�K�,��xJ�֟�������0[Z�y�|B�@勨���,��1.tL �	���mz�

�r�\3�wq�2ΘH���I�F��q9{��b`dL&��WS)�W��[�����6�=䮪�ٕ�"����1!5S�������X�����J_�ZE�
���a�I��7�G0��-b��N[}�w�&��x�l�y-Y�i�Hq-��=?:zF�Hw4�rFφ&���gC�(h�^^��"�O|>q� \*��-�鱟�ó0���nWO��c .��/
V��7Ʋ��@��ys6O7�n,���n�,�m$����������,��e;�oN�y�eۣ�t6�A�<��[�725���S$� I�袬�3�ܫ�t�^S�W�(|�5��]�4H\)���ɑ:0���U.�aTC���s�R}C%�������ږ�dTl6�%o\�]�y�cì�fL����/��c�[��4O�\�#�e~�9`�vK�yza�dk>G�<�W�P�`Ir�'�]a����"��=e�UA9e~p��<Xye�2�2V�o����ȕO���1�׆uΑ�6	�h��ZҮNew��F�g�n4��j��J(-���F��2	4dZ��[y:..)Q1RZ�5�� �>Oew���3�o��G<���"����bRX^���`r���Bh�K�.>�-U�pڟ9����N��4k�����}[��+d�}*/����)��{]��l,J/LȦ+b�q��nQY�O^���Bc"�8q�K'jQr�K����f4��D���V.=��AU��=e�Pى	�!Eմz�����#~Ț!�b\�6��|�
�h�4{ҽ�c����$>H�q�"��.�OW�����:����"�Ox7�b;���p)
�$��K��6he����S��n��Ӑ��d܊�4�L+������vd����J{$H<��P�1��@�&������#���}�MXg�����)-�W,>G.9�Fc�<�D�w%������sTӿĭOL����j�\;�����ɁcF�]��/��Ru�F�ul��7ׁ��w�� Se�b2;W�n:D��'�ie�ٳͣ�R�n�$���م���-,xwȊ	�\'���t���w�����=�O�IQ'�ȃ�m̪ѿ�C,?���_k9?��%�Zf
��Q�ah}��_�挓~�]���o�t��S�~����f�l�ȷ���d�z���Y�X}f�O�߰��(�w�k���-D܅wB��Ewy������Fw��{�w�WXJ�Ur��T*x83�v�V�T�$�{o-����_��iƆ��:k2�j�`�J�3Vv��y�:\�6�h!�G�D�����v�Mo�,�q�W�^٥B���N/���$l���4�b��!��(뿙x~��JÃ��ǖ����S��Ix��/D.C�x��7h����5��6`��@"��/^u��������ב@�aϏ/Ls�y���:������?;W0�Gu��ǔz˄�]w^�K_<km��7�S��W�.E�&�x$~�?l�L��x�-K��O��������Ի��<��򅃭�q�a�B���a㰃�2г!�	io�����ζ���� ;��%�@��kqR^�F�~J���3脠|��u���L`�Ќ��E���X�  �3����ke��d����˱pd~�עh�n.Ń�F�!{�\�{ֱ�_�x��y�}�������O::U�$�ݣ Q�@�P�A{�ss��b,N��&���♥f���;}�ӻv }}5z���»Ԁ0R�/ڀNa� ���e�]R��E��5p�.$�����i��h�U�|��yL@� 	��&��e�I�	>B�I���Q݀����
�M�=����m6����`q�R�)����%r,�} S7�;������]_�}�P���� �d������W����N��a/C��P&�)�� 1�Հ
���T#E���&=:�����;���j���mkj��NR�J����� ���$�'=	h-���<z��M��ђh�A�L��ħ)� �	9{s ��/`���Q���٧�Cþ�Ϡ��.�fg���p���ДC��fE6��Ufk2z��KhD+���=�ʱHٸ1;gA���%��l���יgZ�n�كP*0�u������EM����:�vdt�f\�c���$��vNP��(yx��������%'���
ɒe����Ri�	�#�͢$p����Y*ܻ�'���٭�i�]o�Q���7��P.pn��q�Mf���.�<���P �F ����/� ñ��� 
�D�/F��Wg�Z�ן��I+T|Y�Z`����9���gXg��N�#��Ra�d��Z$,�8��b^��*'���o0i�ҝo�]Fk�ћ�EN������A��%�n�]����2z�\_H�st$�k�A"y��׻ b@<M+\#��q�m��?3���#�H���<KFH���E�\��r��W�4�U.� N�4�R亟"}�8,Co5F�Ss�p��nh�Xr�*����?ZwA<AN0V���^'�l�QD���ȱ�ɞ���v5�j�V�̎Ȯv�d�;KƆ����O����#h�B�ƍ9�>̔j2�%��Ȑu@a=��$��� ��.��s3�%X_���W�q��:X�>+�%�Du��-��a��鬴�j�7oo	w����F�4����2�o� a��3�ljV��A,����DH�hc+߸!�9��@� ��V��|�w�`&����pJ|�hO�l�iɞ#��s�PA�R����mer�&�!cC��Y �\��"�&��f����A���#��ݞެ��^a��R|u%��É<�݌�(+LKQ�p���H����#|���M���z�B_Ie��+�*<*c{�"(�ч�@��D���gexsśT��`/t�Ϊ͢�x��b֨���t� 1q��M�o���{>�9m��w)�=�PUI]m�#ht(�L_���2�QKJq�S*����Nm���]�z���=��;��+mf�����`�a7W��ӕ	L�[�+L�$�&�m)�q�c�'���Oc�%ʸ��
���\��\p�D���'���#~���!F����(��MM�Nx��Eĩ���6R��+Us�/���Ǔa������K�� \@Z�u���8�w�u񪤬ͨu�E7��I��i\��]�r���71:c��Sa�n2X� F�Y��Ƅ(m�Ӑ�O:ݷ%5Z�\�r��-���N�x�0�=�Si�]�
E^��O[X���'�meCZ�X�ϡ��4��Ɵ(��&�c�W/V�H���	ʧ��F�Ss`� } >K�JN#��7C�mM�o�Ȭ�~�r�~6
n�hQAC��=ۗ��T��g��,�
�"��?��R'e	�iմ��F��F�+��R�� �F�s)���ָ��qZ񀀁]o���'�5ũ�p�U�IB��h�(Au�'F�S#���|0d�-)���lo_��Aݨ�\KX�{Q!�Q%�����$)F��f�5�eɥ8�!��i�-�²t�~uBs	 =B]�7��K�
 D� �\� �F�^�lK٥�m�Ju��+�5��� �3�D��ސ!�~s������ŷS�9�I����iO�8�}2��b�N��_s�bR����{��I��6�[OZS��W4��y[bq>�8+�C�������-��)(��P��x�ږ�9|��K�|g�+��	�:_���k����ʨ��e����l�x�:1KD�t6��t������"�2����f�D&�R�Tq���Ȱ彂͑G8�0�_>&; ���n���ɚ>��$O8W�=b-RI�hY�(i^@��J��ԟV��������\a��B�eˤ*z�w1��4�hͨ�X���:���b���d�y��^�����^���m��!�CQb��x�J*��4v�Aēt�s�o�D��U��N���- Rܮ~�T�z��P^��p���6�*r�N�h�����<���~�V�	����T��tkb{��4�m��i�C4PN�9�a�ѥu��=2��|s�\fjE�+��NД052)FE�ܥ��x4m/��P9ڇ�c�8:֖7ثs�JI��F@3��hH�	9�}U�ZK_Е�Q�d���?���	�IV�"�@5Q=�*h���3W���z��C���i��J�Y6ũ����&Hc�>���w�A*�˅�ǉM%�n`�`��_>dŲ��`��`��^x�R������]D�������g��-p�>����ɽ(�Q�^���Z���f���qh���t�O����c=>ja�j����&I,����9�����qèҦ�+D��'#h�~�õ�z��Q�M0=K��CH��S�&Hl��6�q��T��ǳ���D\=ѻ�*Ҷ�Ț�dY2�T�m9��/	t$*`�V���'@���f�9��^���ҪHIn��)h�a�{�e�eh'X���\-��%��DE8JK�LXV2��]C_y�=�|�XP�"�������ֺ��g)�(��@V.���6��~VF��X#E:������m��c|��r"�3��[�>JokV����z����@�'�ŷ���j�!�Ve�]C���v7��0�G�+� �"Fx,�oa�;4�C�ᯁ�c)�bi�G�ҶJ��^�Ny��!�Y��_,��V�3�R���%��j�2��r��{Bm3���t�����5�KUju�>2d��wB��	KH��B;�LS�>�|)�,q�ˉ��|���ԊJ.k1J���aDm}�D�l�/���aJ@���J�{��M7.�1�9��`*�-��T�t�%�Xd����֝��Z�8oW���f�t�8�!XjBb��O���^��&��X쪯����zr������w��F�/~�s��cU1�K'l�8��5� �Z�����Ҝ��g���Q�єe(�����w��嶧1_KM�:���˾�V�����"�٘�Gn�nZ���?1��Ip�JV=c�׶h+6ȕF�O���4̏��#7p�"�8����h�_�&"Uƥ����~�E�'[�L�Ң��� fu�_��������Nac�[��l�+@$��9�z���4�"i�ݟZ兩�^%�[1!�Uqu�����]�3��:@���e3� ���0�	"7�]^CFc�O�8��T��KZ�R�N�F�@����~�Fb,�%�����ʹ�b,��t��']�E�����#n��mGF�9-�bt��k"t4�>�u�L�{���ӭ�v��A��S�>���gښ�KwZl�	0�������v���/�r�P�
�[U����q�4��l���*�.5Ƹ��M��xѱ�F:U�.1:�XF�[Q��!�CH����X�	�����\�oN�t�,�	3�I8���������?m�QF�PW�^��ڼS��Q����D�HfA�}.?@GP^����VE�����py�H���8�}�M��Fv	b��� >닎���(���y��~Xl
�|(�Q�Ki�#N�&��`s�I��Dv���õ:T{�5,��˟{�� V@̓��}���҄Ի>���{^QΘP2E<��*�	�	�������]Ds�\'���Br^ݓ�Ǟ�y{�vEd���I��%����IY���`܅a1��.��+�-�b%]�/7S�v��Ź����*W�眏~j�'�^�%��lR�==!rH�Rʉ&�y������r�0E��]�|Ծ�����;���Yāy��[!��s�?p�L��7��hBL�Pxz�Z
*���u�qo�&����2e���kNs�;���콯G�����%���$���0
ޕM��W�Z��o]�(���9���091]i07�q��y`Y-hf&ނ�V�y5����y$s1]��c�NR!k��{ҍ�1��� �Y�X�^�w���:�o����ӵ��3����o��F�o��N\T뽩���x4Ҝ��R���d>b��W@��� ��u�j��x R�q=q+1]am��(鹾�V��jiuSA��
M���g�!����o���ݐ����<�"]i��-��/Y��=�g� �P����a!���Y���FvS�a�K$���L D�B*"� G45Yw�L��ra�;��={h�Md4|smoc���]����7�$��.r�V��`��%2���e�?È}mP��A7x�j�� ��O ��%�0o�u��sZ{�+�L�6,>�S[cq{�3L�? M���ZI�gS>O����07$�����Åm�ң.�9"E�j��ͥ���=6��&����Oeǌ?���b�;���+���nsc&.S�l�(��Rn������Lc����r�c��M�;x����?�$_>6>.H��u��(��h�Ge�Y���$~:�lNKki�AUK�澴If���	%��Q�Kâi�U�S���� �{*����TD�ˊ|/����0b�f�P37T
�����td��Lj�!����)Kg�>��( >5��FS�����J@��aI:��jg���˥��(� �Q�� ~���Uu,��� �dEl>V�t��ft�D��G�$Ca8�!@�*��B'̂�q<C�em^
�B��|P��Wx����gU�v��9�
KP�3@el�r�_�y���"���ߝ�h�m5�H�Ht���3FG��Q���W77�u��:�O��i�T�4�'�B��T������p��,�vRm���]��OL���]IQk��i	��5�iV�4y_����<�[Д����I)�t�����8H�<[��Q��r�1�+Ue���1�Q�X���<I){��w���/i��3+���}��Q������5~r �؝�~�9���Hǽ��T�ԦU�B��VD���N.����;A8�M���ڞ �D����0	�ua��#h��"�Z�~���
hVٚ����c��#���� k��� ��5+�3��k?��[�.��JJ�B6�<|�����?��B�e¢zL_!�bU���8K���{�o}���#�T��5K�G��,G9�-`��!2�齷�if��!4��tB��p��x��{c�E��;-_ud�[��q9`�6ZV�s`T1��h��u/�貞�#���#�c�I��w"�f*L�c�Ō"�Rf饿�|$98��?��{"�tY���9���S�� {ض�(��z{h� ��װK�U牙�̋�-	)��߻l9����ΆntOK|��ɂ��o�	��D��>x�%�"��ɾs2��ԑ����ys��#G�����8�UN>�lzOt�H�jF��"�����gQ�vV�F���n�5S�;KD�4�(S6(V`)6�~��Gz�����9�鷺��>=�3u�f���%Ȱa�7�����"��1>W<tq0xӌ���B"��a�C,+�[��/��_I�]�kY�(�|������I�>�\M*��w�>a��=�d)�&�YH��eԳ�z:L�����rL��B�a*�gq�7���Ge�\��G����.�ZӍ�U��|&M6�� �����J�{�G�WD���P4�oy�s|k��>;3�ܩ[�V]�#կ�jD�W2��6��3X�7d��Z�C��R����g �.y�\yp���K=8_�N�\R�:[�A0��߃����}\_Z/��\Mo#,$��+J�����n'���l|���2�$(J]�x�L@�n�E2�d{zv�԰An�L#l�Pz�uh�"*}��������H�pH�6��٤; �*�h�"�r����3�8�-�0�?x?k�Y`�E��=�;��j�id�.)7�T�[�[���f~ш
�;�0o���(�FZ�Gppr
Ѳ�s��Z���W��ۨr��	p�+��P��梕�Y�&��>����]��x��[NDz{���"xħHoZU\Q�
�}��B���w�s�x\�b��+�I]88��J����'��JQWP����������w�_�g�ug���V�f�ڒA�����Ӎ��>�l�+����j�H�O���N�+Or�)%���î@9�074w]*'��t�'��D��V���(x�� �.���]�C􎿭�ޜG2���M @ö�r)�"�5���Ьr]M*�I�9+��b����[��l:���7� ����K�'
@�o;]�]���a��_��±��|��4����Z���&��2f�.�F��i�r���y�9��0{��Z��90n]ȣ��I��P^�S��mG��/��I�.��Gl�tu���-��d���`nt!8��r���̬�W��߀y�a�#O'�<hMf*r����<ZW����٢��T����b���	k4�C��#����k�m���,՞����j�����Cܼid~f�X�qi�5;]�*.�>~u�~ll�oy)�=K*���7mA�2'�Ӷ8c�s2�A�a�N�i�e���1@���������&dC���&��$���P.��K�q^	��)T�p,,
� ru��5�Z�7���J$rz�{�B���t/��w+ϕ]�Aҙ�s��B�����oWD*"5K�"�ޅ�l�c�*�ZTI�+�5�U�*�2A ��ۗ,��5/;y�j_�<w�a5��gg��u��m�/l����nl���@;����|��P'�ݤ_^�ʛ��;f2���P~��6�!уի����2Vr.{M.�:��C?���Z�W�r�.J>!�B��/@o���ԙ�^��H���&R~x-��_�Sv}`6]����RHC�`MP��?��p�1Ż�0�@;k����84��	vaNV�3"뵺�^�I;�q�o���L��#�}'�GΚby���f����L�V[���x|�b�܃�=�w}x}\R��������6(��Na�䆷xsA��:���s��-��V�I��`��u(@_v4�7E|�E�.�G��ሶ�ڻ�p�s�[�����/PdF��rLkV�m��AP�A> �}������sF���|ϓ� kO )��r?�B�>貈�D��'�F�_ȼ�P�O`yP�`��::��'"H(�)IQ�;n��WCy��MM���9B5�I�sn"�S_�QX$�z
�}���(�9=�'�[��yq+�b�M�fa���o(�?�`��%����C�Z��)NGK���}I�Ā��|Mi�׎�Ļ�M�Ǥ�*�UP���i�̠�Ӹj;QV���Hsp�/�^@��Rk*��'�Q]"~�B���"�&n�m? ?qG��H֊��_�W]� �(7�D�mk5�ț4[�1�E,�03WOt2�b�
�/1�-��dZ�[5����w7F]S�(ֳN�����&-
�1^�$]�G��:�G΃hf�_���f�%.�������PR]��'� w������WrߦeT>��ڪ��΀���h��ڇݏ���f�O;�쌘��V�$e<B�#��!Ki�-+�òѼ��	/i?�����X��o�4������L"´����� Wv��1��XE]�ƞ�^];2�
{"��k�8 ��!Ş*�`7Rz�U��n��ز�j&�E��DA�gV�a��4�n��2ױ��
��C����9�$��	juf��đ�D��m�[�%��8j:���Y�6�ns�.��-,��n�Ў��qf��ו;&r�)\�Z�Ú���ak��U�'0�t�剻,0��&��&\Gt7�<�?���md- `�@���Q?��_Q�;S�� ���� �7[�LPp.r)N!�R���Ԯ϶�-i��O�ȼ�O;CJYY��(��`�=pԹ5�S�SR^�����t�D�1Q�>wE`Q��. C�Z����HE�C#Y�90CK_SF�$���g��!��{]697��.�>�g�42���<j4��Fh9j��c$稳N�G�`^�"`Q��(����v�����H	�yC�x�s��b���CݓP�����/�@���v��ż�6|$8ΐbe�j�g,� �����+�S�r�l�
�ez��hՒ�+�3���ma�ٺ����-i��Z�O��1ȏ�fo���+~A�m��3`�g�W��ixצ�ٟ�/��vJ`��O�'p��PD�eۇ��C����<�)�+,��]�n;#�/�@�Eb1����AA8�m��_�Z�����%����m\�ݛ
^WZ�j��4��Պb-�cx�Q��VDMEL�pF��� �����x�5k�Um�5�L���合��YdG���u}U��+=��2��/���8���L����cZ�{�jA �ݡ�ͽq�2���D�sA�����Z*j�b|�r��t7f+�$DG��DUfN�[Ɔ�B'�,�,݋�����
�u0i�g���|�9�w-0�a���0�n13#S��W��lUv��U��	?y�猖��G̃,���Bd"�M0�E�
����[�e�M�us�}F�H�f��ל��.�fkР�c��B��6�DBDJ����#o^	&~�ِ��`+�o�c�X�o1#cG�Rι�������q]@���l���#N�D�3�{�A���;�8����/,Lh�Y�R�(�:Dl�΅��g�ƴ�x�%B�1��%�u���c�/^�(�7�Էnq��^�D���O,LݼKa#�n:��P���$�;�94)>g:tAiL*"��5NY�{C+#�`�^�1��ޣ����S��Wp�!A��?��d��в
=K9-��|_�;N�Dl9r��{���g��*����f;�N5%�0!���$��d=����5�,N�1���f�����IF�aa�`
����U��n�&�!Nh�ߊ�ICo}�6nJ��è�A�ʜYxNfd��,.�X�^%����0~ĹpJ��Δa�ot��+_�1+�Α��=^E�ud/��e���Rޮd/�s2� |5$������e��dtZ�"��{zO��Ds��ƻ0-����XW�'*�7��7�V�[��o�c�j;ӣ8T�H!t�v�����6=އ�R��cf����Z�)�tv`Zl�TN�H���4����3x�2�6�L�8}�rF�*^K��qtl����=_�G�F[N�4^�������|)mL�w���0�����-���D�����.�8�
�LJ�{���_�A��oho����M�$��pK�>�~J�褐��$ب�oF0�jNDF�b<�=1�#��6��ת�7�;]��Ā��R�a2�Pہ�B1*g�V��>����J�*�^s�-��_�?��.'�aZDf<�qJ�(_�t�w�"��Aˀ�����9���`[ydFu(�BS�QY5]7U�(#�=�vߊ"z��}�у�EDLU�y��²d>h3�"�0*��W�WI��~o#�j��Zc�xK�h=ܧ ��+����}��'>�&��hvW���}����E���I��ϒ�.I!�^��"��<`�T:����V���_l���b;_*��exi�Qc��
���f�;�竳��g0(�|k����*1U~&�����ԅ{eJ����"����#���������=�¨y/�8m�9�5�r��Ѯ%Z8�kd�a!�������,�{�UH��1�\��;��W �<l2_�IĲvL�6<EL�_��]x���"c��z\��g�N�P��b��J�����7	��G�2QՅ����7STgϔ>D��?�p��޻�Bo��,/
řW��܊�����,�,@ʐ-�����!���3�a/U8��FC����:�p���2"�:ݎ铠#����Mz�y�%������y�1ĥnL�QU]`�5z*1�jL��0`��\�*!�����2y���D.�)M	�x� �I^Y���"Jl�W�
�W�J�qCp�$�6{��5��;G���f�3}�IhZ�Nk��E*.��(%���ݺ,Z���\X���nP��b�����W=���t*��p�^��1���4�(���&��{D5�X`"��l�J Dc�|04t��X,�?��`��w��#p�����#^�W�5]�&��9�^ 0�m� �	K7E�D �f:��+ם�)�yqq�׃��;���ğ(Ph8��,ts�@&`���9��dM�R�P�˞}��Z��zsP�m�Һ�Ƞ����_�xǿ��].i���<����Z/͸o�'�pG�ٞ�Ζ�5��ϯV(���fo]Piٔ4V��I͟F����}Ëԉ#��%p��i�E����]��<%"�
&�Cu%�j7�0��
p�4�c���_?_K�E]T�]}�U��1@�X�Y�%�ΨkBA=o��[#�X-і{��- �~�L�M-�}|
w�}�~�Ŗ?a�.�e7��R��Z��?\�0�"ڂ�Վ^�ɡ��mu�"�>�R�Xl�,muӘb�Sڑ:s74K4�� }M�'�ua�B��N6�?��v�;�b���g�?�
O��=f�l(�j�����fܱ�N's�f���8Z��hz�d���ZAL��yz�E���[�v �ߪӝ�q���1����Q���W����t���Wi�Ը�o*�v�q)�S��Wo.�61K*s�1"��
(�蘑���$s���X��XX�v@��������AJ���U�]y��H [X��-2	�~���g���4m�%L
�������wr%��&���}��0�|�R)�k�E�9w_��yu�|��/.:���*��.��pEv�'.��B�DЇ����x^�c��j!�-PJ�o;�^����5$��~Ř�������F~ 45� d�r;R�*I��%���G��Q���������^�}#t�&�f\��t_�$�kw	2}��:���m;�*�|[����9=��V��JG[< �����<�Q�1r�ם<"ȝ�$��O��E�L�`��R�[;�Zܗͽ��au�t#E�ڊ�2C���~�ba��L�O&d�^1V�OΓD�0L�9��:Cy��׆��	)��Sg��#i��!#����@���Ek1W/��k�$�X�χ�HiN�@:&F������5�G�����T,J+��T��	rJ�]Du�n	�3�����MQ/�A�G�v=V��T�ʓ� ���Vce��̊�);���Ě��oz7O���1#��;�TI�в��z�H����د���a�n�έY���,�����i�hQE�J�)ѿA�L��^3�7 ��9t��a�F�6��\&w���(�m/���ǀri7�ʊ�F���%S`��ʑ��R�{�}G�%cr��Jo��p���$���tK]�t�k��Fw�K�R�_�t�N��e�@�"
+^����y\ߥ���Lp��<M��/���.��d����% �X�R3���	R7���5�#HIE��v������m4��2pЦ�Ց�E� �
�l,���j�>k�\FQ�O�ȍk�`}��3��"`��b��&�A�B��G/*��&� �~�:t�> /��ragz7!Rե<s�as#�T��!N�s,����#�ղ��kk��L�e������%-�|R�3#,��	���Zl���R��[��#c�9܃��c�w4���d�K������yW�Zw��w����y��M{C�W�3g���������O��̲̀:���c�u��/-"�Y��hO?,���}����Ĉ�&̍"<�LU)*i��V�2y�q�1o��ۭw'v��r���NmLPO��N�#�G\C=���:5�-�d;>��OQ6���Y�c\�C����"�������3��ww�6e}I*������L_�P�O_�����R i�+=�yi��d��.]2����x��y�C�|�fc�Q�ʲK�'p�ֱ��������T0�ޒ��y�;,�{}A"�4� �l��~B�Rj^'u�J&uCG��Z�[�#F���L ����Y�vr�S�J���9���n��%����y��&�����ѐ�2!��1(d��G9�%�8���Q��2Re�����E�QF2Dh��=vã	����Z�iA����h
p�P� �]�C�ԏ$���{�P9@��惃F�i,�L�����[��t�a�����)!�+��]$/Nlt��8��E��閭N�hE�1�u5�]J�.e��n�l���O�V5;i=���rǊ�j��Dl,p��Gׂ0������F<�hKA���+ί����;C�e���2�$r��\�Wʇo�}l�"�|DH�)o�j���x�S�9�3I�ܘ��� j�}��_O]]�b;(�	s c�7�d�Z�k>�}����y�niM��a�+�Ȑ.�jX��R�����J>�)+]�?��ćS���F�V!�����<8�M�J�wb-*�+�����˒X��zz�_l�H���U���2^���ߓ���F��-�'ҥ�� jϴ���f�<����\���Vf�ƦR.����I����-d$�iC��cTN5�I�g
���iC��,��CZ1�$Ζ`^<�Fp�,��}�b��FS��;X���eH���fڂ�?,�{�����̄�j�_�.��	����g�I�v���3q1�潴�N��"��Fkk�</����O�N/�z*�g��,��=X��
�fĿ#-0V�rb7��CE�\YR�qK�W��z����i������ԯ�ƌ!��>�C�����7�Uη�	1�W|L�����{���l.UG�#� �{�t	V@���l��� D�~?u�]�9��<����q�=s��h ���;?�S�i���N�/�o7����k?֋��	!�Z�o�cpؽf^�_.r6!T.k��y�ɞƻ��ٳi���e�S�z����U�#/M��������ҒP�^�/�z.`Hm(�N�e������)�Ix�ƷЋ~�æ�Jփ�O?�Y�UQI��� ck�-$6����+ô�	�ܦE���@3J�mn�Qӯe��LC*u[�h;���C�^�|��^1��������~��e�(F��uX8%�Z~��P��P���ꑯ��87�*|�H�}�A���C�����Nc?ҒP(����	�Y�f�e2����
`�%����F�a߲���l���ԧ�lE� ���#���σ�k�,�V�׮ԩ1T%���� p�q�)�����3P�Ц���߾g�հ6�F���:���f�GkKX��5]�W�W������c��'�K�uXR�2ޠ��0pf"pW��D�9��n�u���}P<���W�&����ܭӳh�l0~�!i�=s���	q����N?�O�#�`<�,2���,;�K������ɍ���<�<��M*�����ο�s�r�#&KYyLhw�t���~��?7d汗�ǀ�ҘAhdh�z���G�[|��Q��xB�5�W� ���J��1W�#(�v�����	�*CKQ��{E�780�_�XvO~ͲĮ�B���a�{'��o�VS;��Yܞ��d�z�_19����"ފe%���앏hل.��r�&�����b��X/V��.�H��n��w���;be���/�*w�Tk��W.��s?����q���D�`>Q����pq��I�$l�k�.讎��ˀ���U1�SX��Q�U2O	���{&_>YU6Zen�?�BU
R1:��0��m���u�e(N^��R�@S@�����G��>R8�~��-�P!cq���^r^�	䈎�귄RO"J�GS���3N#1�.d�l��(�P�9[��=��dNБh���+8�U� e���Zv@����P=����=J,���<.�y�7`eF5-�d��?+ki~O�?���=��6�cWo�;�u���Rn�O�7��I�ys&��j����-u�X���U1xl�(h<�=Ν9{L���5◂)]=i�]�ez`����r#�3uS)���L;�a֤���5lh��&9Y�.c+�G�4�8�3�Ъ/]_�)m�F[�jv����k(��lV,F`�dJ������2!��jy>YȽ?�d'_}F�� �}�D�Ir�7T���Յޞ`���+j��E�	��?v���c��q���no��Zb��+�fD��,Sd����>t��IZԴJ�����iz������,�U������1���K4]s�Fĝbaw{*��N�ȳ��>�f �r]���M�,���m�H�=OX'�[,�g0%��rTgƊ%�K"ء�t[[GE'��Ť�@8܇`���g�h�Ҍ��Hħ$'�]a�f7�S������@G�Hc0�k\�����Ȣ�#����m�y~��+!p�̳��H!F� L�ʟdS_坫�q��h}Q�5WiOߵ�oJ35
���K�ڲQ�<S��Q��Z��
�H����Y��MI�ܸ�V@��ƽ�2"M_���21�֤������h<�> �D�1hd�Rvf��Ϝ�V]�Q��+����;�����*5�lހ��>��-\�����p~'P�[�O�y��zǓ�n�Rަm��vo�{�=1v"j�w]�:YA|I��} �����8Na���W�\2�x� s8ҩ) w���A��Nq[?J�%��ۻI�1���oW������hZW]����e��b�����Zgs�f���Z(��IQ�2J���r��f8�3Z�
���Ra�����sX�`N1�� xJ�L�z�Ă���)�)��i�e˝�k�~��ߞ��� ����+H�8���������Zk�CS���mX��V`��
�^9��S�[m�b,z��9Im�����s���́�8��	G�b^0��;����(�:Q^�+��}y��I�����s�$f��_=�!c�C��F_
<{���ێ���[���p4���!� v8�B_OaNڂ�����|q�~uS�d��\;�7�B.ߒ�=ֳ:}�|�5�*t{�Z�V\˼Ǐ�*�H$_�ɹ�,?^Jګ������axV���MG�zz^Ө������ո�
��M�Wl��0
"Z2��E�}���R��ٰ5~��
�L��W-�2��4�ߖ���zU����޸*�X%=f�P�����|���P�R �y'ki�Ձ���Br�c���f�=E�2>��;R!^`Z,����@�*�յ��K��Xd����(W�a.�k˔���t5�	��B�nG�hW�jn�3�={��w��4GH����x�UF��h����ާ����ښc:MeE�\�(���}^�����g��`��[�Җ��W?џ�lx�vk�FjJ�_	]��O)ƗR��3`O$UJ	9���Z{3�8y���]>�	��50���%���G'P�2��:�v_��oKFJDb��fmH���T/H ��A�$�Yw]=����/�Y%��;y�M<>;_-������%7���Dk��wt0��μ�=,�)�vb᜼e-՗��WjDz+U�?�ؤ����Y�]�����
K@7������@N��h��
:�r�F
#aQ�`�C{�=���_�0���`��"��su���L����,<F�l��� 2w���_�j�Ο�B�=����mx���!5�w(��׺�ɉ�ӣ0�l@iCQX�zb�3l� ��7��t��������Y���a��-�l�W:��|��׮+|�,�Ї/�>)%�==��F�+����nl�*����y�o��(R�mD
� �S������x����`��"?Ú@q
@�Ⱥ���(Bȱ9:G!��D��<[󯵾��z�1j��9/�$p;����ĿB\��XJ�BT!Ҭ�{z��=s�<D�Xs��4s����[�#O��i �n�������F���e��>�i�0�`u�C�$�.��G~���
�����nҢRd��-K@��-��Dc
�#@����I�T�8x;4��,\x�!rbŬ�3F�n\�}�19�C�';���?wA%�ύ����r7�W'z��j)~�B�[�M)�8Y[s��m��W`w�>��^F_#^�I{Z+X2C�� �	A6a=�°nqFM|&�������Q�}��r��c�����F-�����_�?��gԽb�k� ~��:S'�T	�ѯ���i��
��[	�!^��h�
��
0ٱ�	&SW*��'m�5 ���K�V`��\��&��W���}�&��V��dr��\G���0�����bu��Ü�=(�bYGV� �y�0����J�$��`E߸	�|�n�S��%��t�na��|�*>�8%��:�n���g��ҭQ���#��i&`J�d��@@�
��^`�b,<�m���nu�p�Y�]��3��(|7J�aI/0G�I�C���zd ۼd�����UIO�ўR��|����wRv��jcU��՟KR��t�rV(Q��z�f�25|�>�腦V����};�^I-Yj'��M-SC�/E�Br�o�V�����=LR`�f�'F�z�� ���R�3T����#�hA��ǚu��mF��8�~@<��}��V�m΁�f��}􋹻`ܣ@	�ǅ�o�g����\��)�G�E/|n���c��S����.s���E<mlG��6����Vr���*�ޟ�� �Yh�T�Y��Af�.��^�@'�h���u%�|q%;�F��I�J�\���d
#R-9H��ך��j����f�������
��_����JԿ#�f�J5؝��lߓ�� ��ے}�� �E��2�r'x��Lo��`�`��F��@8V�|/ñvx�T�/Z��Jn��Y���"��`���.QR>JM2y9�|Ns=��֨�M��s�#t|�N�7tj6��YJ5K��,=H�-Iɠ�Z(�F��,lԳ\��7 \�)Fy�Ƌ��S&D���PT�{�Y3b��	�O4����?���@b�]ȯ�f�B�t�����3:��f�ӅP��w��0u<����Ǭ0��d�����6�����)0��A����PA�Z^��ʛ����A2i3_z��Z:\���A�䁔W#��x�W�I�q���яܘ�zg�J�Su�<	ɢ�P.�u^W�q帣iy,� :D���V���.HG�����rnVzA����,���M46<�y��ݸM"9u��q��D�f�yiP\��|�x+�QY�i���N�N�����M��^�)�%�{`���[*N&!�*�̪�	����9��挞�x��*A4H	 E]k����s��Փe��^}�`y]t\�6-��#�7+F�&6��x�uy��q%��26&9�:��!�x�/(Xɕc�.�O^;��;��l����F�W`���M	e*��ŷ�*c�If@R�r�,�`)����F���r�Kptt�ZM��fTr�м�K���L�w�^�w���g����&\��vl�J��OC�1��&h���M�-�C�����&�+
[�jU6K���&s��~c����p%$�J���]��V3��<�m�QCaZ���i��!�zW|7�ī")]�����@%R��e-�n���籺�{"C�b+~�����G���6�%X��E�n���̤�񯭧d�0�G��**�*e�p,��� ��d �����m]?�0J!vF��1^xr��s�G-���ew˩�G�����{_2�2Q����G�W��V�v�$b�$�N�����l(o����8�@����:s���  �x��c���1�c��AD��"�%�e�XYkk[��#,��ig��E��S@(����ʛ���} "s/�'��z�z놇�~�=a[���x%J�1��ŉ��-^��I����V�� �h���$��J#f��cr(E�B�
��No��g��bŁdf���G��-���=�Q���J�]*��.i������(�������B �<�Q�j��� ��e�zc4˓|(�� �%���5�r��/�tN�����p��5�9�e@���+;��<9�� ����Gbw�;����h�t��)��u}�q��g�Op{;ɣ'�w�d+d���}8�C�v5pkc/������ܛ����"��NB�Uӂ��i�n�V������T�u�u}fFf�Y˻s�,�'�7#0rH<�Ŀ�R��SnNP:��9�ߖ��M�;ʦC�һ�o�h�(����������+1��O�8�&J�p�-�8`�)d�E@�I7�F=o�7j8�%�V���}��?�y'�-z�Ġ�.�I�;����~f��#�_��6&'��ޛ����k'mӢ�2m3�v�km픈p!�l��&~;c���pm�*����Y�M���RX��m��\4�s�BN8�tU0%M]�&�L���A�<R��B5xZ	1Z�,
Rl����t�����������_�IH�S?�Y�t���K�����P��|'D&2�I�ˀhGЩ�y����O������m�2
�@Ķ����o�J8E�]�N��x��:�7�ͱ;�ʤ�*�V��(�2����'v��/��@	�¯��V~��;n�p#���N:n [J̗���XN�L�.�h~�?/�A����i�������q�i�;��'ND�U�������я�>>,gtQ�T����&(
�b��_��}(�O�HW�mr����-�+G�*˄9e5]������#��ﾨ6�,�?���FP䦸�1��§T���p� ư0Yk��zNa�o��K��{zrX7��^��-�jV�GX<JV�!�F�n��꿅h[2~\A�Pv�/EB��eh�Q��
8�p�"Etz��8ղ
�5��|�|�X�2��4&��Z���p`����>I帬Mq	��S�cy�K�YJFy��8dm�L���8�f�q��Kaj��'C
�Yxu�Bw�Jp�Q��+k�Î�����pu��7Ѿ(�OPmzxr�� A~os[��;�%H���BQWꊵ��o�U��]
��X����P�H0��s2@�g���X|�s�\���&B��H��Z�!���L���L�����74NA�j��>���F�J������U`����mpw@���2�+���#��ڤ_bF�Et�G汯���JY��6G6B�7���f�_��I6�=�AL� �P���������˨N"ޕ�� {-����SdwSY�i�4wиe\��G�.�	e�>'TK�1�w�}NZG5y�M6+�e��V�(����귨��UmCp�/��������sE�wJ��Z��iԱ$_���F�E-�_W�[(����d��a!���%%V��|�����	FΠBK��"��sJ:U��-Vʳ�3�~#�6��@�	u�0y���l�F<C� q��,�I�� 1J���Ľ�@���ݍỳ(�ޛ�h��>�tg(�{�mK����+��2�W�˯:w�PP+3j�����2�*��T#�$U��^N��J@U��m"x�IW!�w؞�Zgۇ	]O�ї�q��|{�џ�ít�y}I=̅�	w�z�#���m �DD|$[��`$����?ф��j��C�砹�>yH_��ƺ�5>����
ʸ�������So�P�v�]j�Z?IM�䲳Z��XW#�"��X���
�ʹf�i�� >��	����"눖��b�[���>�	3��sca�t/4�����Y�1�˶����n�'j�|8��_���E"�tf�4�%Fh��VX*ҖE��p��p'v&)��!�k���������tڊ�����<������U&�6�E^�~��?/�e]�I�`/��D�	%t��^0�^�U�F�F��?�U��/K�
R�^�9��&ja�Q3¡��)R}6��LMY4+Mv�w{1's��M���-��4R�?���/+��h��_̴���MGd�V1���w��Y���@�̉�����C6���G��+N6���a&[]:�tM۩/�%*��w1�W����k-��Z����=��0nQ}
�pĹDW�I������4"n�����:]a���_r�\�����+o��2X�p/A���Ch�A��;��q뼅UL����^�P�/ʳ,ݯ|b��aa^B�b:����Co�K_#�uj~_:��};�Ĳ��%��-�R�f�(��3��Q��fC�&Q8��A (������☸Z�J=�P��[]�k�W+�D��y�=�Kd([9��u�t�q��Ҩ7�}��~�� ;��|��G�V>�
������>���_õo2R��{��5������~������[�?��]����O'[�z;_�e��I��OK7huc�2�#Tc�O�\e��\Ft�+y%f�e췔.�/"��S�X;������wuUij'_�.�|G.�w?j���7���U�q��[����8N��}��*�[m��OP-�B2qU�������x�b�~	a�}K�t����04�ڢ}���=a��na6�<�>U�%�Jq6}n�,�V�B����og�,Ѭ�m݅�Mm6�i�X���\g���<i��������m;>fV��
U �F�9������ܼ��*u�:�=���ya�ti�c�]� Z/� K'l��듬�*��	�gЮ�>N~�1�)}�ɶ?Bs�tt�i_q>.�p���[������ ��N�j:g��H�rf_\tA��"��$+�$�@NX=_K�V�����%���-�D;�{Q��ϫ4�	��UĲC�v<���H?���'7?"�}r����ˀW`��3�ܶS�m��?��a!�W;`cm:���=�㙄��w�KVAP��u������+����h��<��苋�lAmT��,S�����t�_$Z�����(VLް|���5�gõ�_쳊���8��LBn���GK��L��d��*�y['K�k�M}w��*I�D���U6ϒ�=Gf��e� ������O����,�DW��>e�H�p�A�UH�c����<*�
X+��h�����D��r�"1$\�IY���]/ m��ֺ�N�q�u�s_�y-��b-��|r��+�}��r�� �
[�1ɮ�S+`d��W���-�8�����?&r	�Qbԗ��삕������<Z�@���X�5uPHݧal�Z�t��=�@>
f�&��� ���Z�W�r�jҌ�bLV�15g>�w���B	fAx=���jh�x	[r0���s^�wVdl7��
]i���:�A�>Vᐓ;�k����ڥ���5�s��4�1ly�����ᒻ�"Kҝq�X�?�m��1��K���v�'�=�(CW6�J����0Q����lP�"b��#��b�,֟�+T�%y,�Q�ߛd�A�؟GOOƇ�@�#��	���*dT=E��6���v���љ�̠���X��'�BL�BRD���o���H�X*b�����0�>�61����!��(~�9��3j�t�y�x��T��>����ɑߙA��/3�0����Y��r�q���+�*\A�e5I�,3�+�d��	��Rx�d+�02�s>��v�/"Uz۝��A/���̾��ִ]FK��sv	���k�/�]k|�T���(m;���@y ��w�hM"��o�=\ߩI�׾�G"n#�n��e(m ���Pk}�Mj2�3I��,��#��f�7*5��iw���Vם�[��Y�{�/��1V���t�&L�Ei=��*֘��P���Z1�ܬ�z�s	�;ɽ�TL#���Ld�I�s�u�f�"-�
Q�sC�2�'��R�H |X�ш6B�R���_EIï�n��&T~�����W���1U�~�B+q�w���g�a+,����e�C1�Do���Sd�i��^R�;����e�U�h�R�u˖���>���%<�qc.��8��uCf�c����Km�f�=��f�W�I^������$���a�� �=[M>ϒ�,�֡(�|���JWX�\�*�"u�!�s�6����W��U�W����7xn�E�Wo��;�:�-95��~go9R�=H��I���1��C ���wj��۷=���N���g����-M�V��!�J� �T��ݫ�(�+� C%� �*�,Z��>%9�wpW3v�Om��c�6m�k�J�e����� >��C��lv�[ψf�W�-� O�㕩Q ��1�;(��+p�N$y#�!�D�0#-s�t�"g`�rR�ҧ�7-4>ux�c�q�y��'�P\�r#CX-���6�i�	��D�����L	��|w�t�w�\E	�mH�Ѭ�Ƽ'P� %}a!#���y����]���9�]�GG��G"�v����ܔ�q�����򃐱�gow�Py�JUB��7�Q��Ԛ�[���s�N�d���9}��PR��D��'�~�cYUs�h_hQ��k����}߁ņz�w���������)�M>�%w,�O��)�i|B,-6�ū���1�w�<���)PU�=����=S����n^�bVYO �yL�R�x"�p�z3Pk��)�2:��&��*�H\�Ûk��M<���W��J��v�L�P�I��̘�qj+s�H�?��`� �o8��?i�[�P<�p:��w�w�\��dN��	��V��p2F���L�8����] ���n��I"e�ڃQ�~�a�=V���O�COz��F�e	�k!mp�4˅.�F�k����,����W�g��X���?�#k:飴���3q4eB0;�]�X��l�'�4������@W����=Y�o8��.�C�$�;KZ��D,���/�}+�ݎM��#\�o��'}k|a���i�wHc&U,���ә"s���ɐǚPX��Q8"�N�F�\+����Xͧ×���_�G�[Hf���`e�Ƀ�e��o�͑+��<���m��2�z1el�_	b �[��'�.�7a\�5�9��X�J7���\Sa6�::�p��9Сj@�6��b�9�co��l�����ܶ(��E��9�߾����+K3X_N��ԄbÊt��3��z򑲺_5v�D$��;V�������Om� F�C�1�� �^Y/��]�[���i�:�Q� �.�P�`�;V������]������-N�Hד��"ͺ���
���ƅP��4��+�����*��kۄ�h#��m½f9��f���%/uh�ȃ�
��Kw�piXt.�Bg�VW�m�~���{��R�(���n�C�$���*<��^@��-�����'�Y�l.u�Ck�r��_��Ãqq�uVP1����e�-R
/�3$�e���i?����>�̡�AJY7��N��� �}��.(Uj9^�tks�c�0ܴs�Un&���C��@�!����C��&b��Y6�J��
5l�� ~[�bvć�B��&���]���.��2ԍ�f�%����]P��g�:�S����V���AyB�\��!����%o~3��.��1�v��q�[��!��\YR�=ٿf��>.&�2��(wf"��\��J���y��
�'��;�)�� �Ay-5���)��
�c_��D&��3�)���nS�U������B|2Y����o��e�O51z���rmM�ɷ��D*¦��>��R�����k���GֻvN�ʢm��B�B���9�0�I�Vv�sئ�Y� �D�08��X.���p��)&8��ܼ��R���j�ƕ���~��i��'7!�I�/2��*hC��F�"�k���M����f���������T_1Rs%����we:���	�B�Կ�t�f��Z@�_�е'/���b�ᖵ`/h�Ğ�Uv�)6�d�ĉ�������F�&1�؎��XQ	{-���vؾƇ~Ae:�	QĘ��L����N ���4C�F��$MβE����~6��M�7f)G�A��$W�-�� V�f�վ�GL����-8��EO��n}��?��(�z�4`Ԛ[�-$)�Acy���L��]9�ҥ�8�58#q�hET�u�����#��Cn'���J��/�c��v��c�m���S]�3�����k���.�Q(�T�]ڶ�$���3��(6� /u��92�r��pI�Jd��ṁ� ��C��2��|��̎1���f@u�1���? ]wS�^-���c:c���
}�e�(}��]\����e��<�l,QW�M�jY��X�٪���&�f�/���W�Z���'H��xX�L�w��EY�|�Cq��/��z�����U��{�B8�!��=�HQZ�&b`(��l���4\�b�a�Z�e]�8�v�r4��"�؎����Om3s'X�?��.�O�7�ȶXQM�7���%%���X����@�=�8Ig?-}�Q����_�X��m�������٨o��#0�����q�����{?RF��%��>����`�5LLA;^�����/Q�iMp�89�/ttX�WJI��ű�-M��r�zВ�;��,	��Ė�"F,�>�-�ϚĽ�Nz��f��$H�\ʻ��
s���i��Y0�BĴr����]��~���	?�-n7pM��qM�w'��(G���9i	F}����Z�3�0Ez#4�?��_�e�∐Zg�l[<m<�$!%�M�2HDJ�v%�!:q������W�2�z�Ϗ�Q�w�	�W��`�찑�ۗ�~�hgK��T�0(ڭƿ�tЌ��aO]�FK]O�)W�ąfKS]
b������F����d�=.~���4�<C�g���ΊP����ɻ�dY::�c��*4=�l�����͋��w�yR�*�9�!x�����v���ȹ[�~����l�?v0��=�J�'QoZ�f�
��T�>j����P�Ͻ�7M������L�8'��\�1ޣ��|ɑx��LGM���+	k� /�TЕ�a=2�WĨ��$%fX<����by�����ۙil8E����U��V>�zd�s���E�%�ǌ�6���y�5��/���y=�>&j����X
�Vʢ��c��	Q0$y�2'7�F�7�����?�1ofT�n��z� 	>����	1$�֍S��d�]�� �ބ=C�{���8#1��im`Cg)�.�ì<U�ɮ�7PAI�����"�\�jL���|�1�"�$��d0+&�}����΅�5�6W�("f1!Dߛ�޿�6���"I;�bw�O�����7��j�P .ojL���,SgSt;�L;-���`���׫������t$�T�Z��c��#/ ���m:�v�"������Ͱ���N��(�c�"�^yЭ�0U�+�����!��)'�^ZN�ktME�;u[�a�_���c���Â��5�&�N_O;e�,DU�ww�_��{��d"�r{Q�H��J��Ō}�/ϴX�Ǹua�H*t�	��
�9
�P����w�W�����`��:�[�4�րeZ�^��t��3��P_z�
p���OҌyt ��F���&x�١O��Uk��]{����I�J*�j�����.~�yXR��A����UB��
�eM��$��_����<�~�1L�oWߨ��k�Ts8��-<��X�8`ROސ4|П�.|�P���.��r�2�s�-��=��L�\��s���)D�ĵ_�MLxڪ��y�5,��-�ՠ�Lb�Q[�V�(=^�����+уcw��A~�V(+N6��W���sjnO]�+�C5`4�]��z��Q��D�q�-�jDTY'e�I1��]��C6/�3�k��\6�ף������^��1�_�e��;�&���ql�/i�Lv:���b��GӢ�~$Eɮ�B�`*0�g���[�7�(����(��z��HF5�*�Su�x-l��Q��k?|���f��ul~���~G����E#k�E ^�,b���#87M?X�+�`���D�ֳC#��mh:�v!�V����B�~ج�8���q�b|��YG�d!~�R�UzƇnn�׏zl�Q_+��@ڒ�l�4�-O�m��jNH>���!���Nb{-�Z	B�M�a���Dɲ-��HP��?mb�S.Cu0g V_�s{x?�a�Ǵӂ��@q�$�O���$����a;�&O��a}`����LԉK�l~9�R��������=�7�{��?��sKh.+��! c���O3��S�3�@���bs\8��mX�����g�>��`�:+q�2��l��ꉶ��; k/�U~��6D�}��ǎX\��}R�=�Cʁ��`�������a[߀_�x퀉�]�_*��B�� G_����'�������E=�%���'�S.;wA5϶���V����A�:�98R�N���5����\l��A�Ymɺ�C��6ȧ����� [m����3��d'���R�0��_ߓ��,�r T�h[��S�H��>M�(E��`Q���*@��X��R]�*G#TH�'��"U;QF�ӭ߾ܜ��s�A$��lż�ι�_fо�Z��	�`>��ay+*/[��`�5Gv��:�t�>�ٗJc����v�V�v�ۃw^࢕�ȏrU�4�5������B�`��/�%�!�_Hm_Qt��Ȅ�}um�����#�'8M��ƺi������|��ƫ�^�s9���E,��E��!��l���J=���"[7e`NwQU��G�؜�叚:��_d�췤ڝ�Qu�_��&��r.�1/L��T<#sI��e�l f����T}�>�E�M^*��l5W�ٕd�Ⱥј��c=	4�d���*��S!R9�=�7D����ܹ�0�qk���\��z���l������pu�D()�����%kPh���M�1�E�
�dSu��C�r�}�<Q��k:��� �Z�5#�,$���@��޽ג�U��X:=3@�}�@9�'7Bl%|у��pGJ�T��x.�:"hOm�-7@��xyn�'��o�
(�E� ~s:�� �K� �^�]�=5M$��a_�&�aO���3���-k��o�MU����P�p��6��ʷ����Cβ�.K�i�n�t�ݧ������G����<:YW���>_�R"W
���Ev=r���ϸz}'�����*�0�ݸ�����O\h�����uJ�{�=�j�ɴ}��~�d�B7�UD#Lk��Y@�1>.���mH�@ �G&|���ZYo���P�`��>���^W��N�#�1i��T�����*G4f�ٙ}�m��/q.�͇RS��o�!-��D�`c�0�����q�����\27�9��'�5�P#,� l�bR__��rs���,���s�fg��t��0֥k�-�ȳ�]'Z��!w+�^ݦ�B)��M�A�����@�\���k��:N� Y��-�Y][O�ؚ�4�T��"ocA�M�xI����X�ԍ��zņb �bn���֣���*&���3-�H{�m��8�iM��\���/��N!i�Z��
I.����ŷ �܀�O��*����>@��Q�A?������S툞��|�z\��K0��\R6
�W�����G�[ps,��\>���ؐ��E�k�͈���y�b�E�s٨֋耼>��c��������\�k9�$%� �5J���?F�#y�|DSP
�cR3?[o�/냫7�� �5z���ث�a�t�B�v��/!a���甌ؙ���d�t�V]�8�O^�FOUU.hx~IBd8ц�s��?N�.��9/]�ǻ�������`�>�EU.���[� ������d�;+�TA*.+���2z��x��Mq�O�8�Z��B@p��/R*w�P� la����o<q����Ϸ��}H޴�ˁ�a��	�Z"O��V��/?�R%^��ܻ.]�G��o��|� $Y��vB�Q����!sYx�v�� D�aO���mIE^1.��/|�W�U�< h,BE>@[�?m��A�`��>5�呱�F�x�xig��(7��{���<7;x�2�}v��V�!]8���S(G�`���3��_�8vT�(b��b){�s�Ygӽ� x�"��!@_p7��w���~)�������5�԰����L��r�+N�3�%_'���G��C��O՞1��q>�Q75�ڧ���(N��vkOv<�7��gZ���>B����J,�1�Tᵮ�>���"o]3V�����E}�w����8����7׿�~\Y|��U3�+��i���7;��fqU�;l��s�~�K�i��+=ďa]��6Y	Yg�K�#p��vt"���&h��5���@��%;0�,�
"B+�����MEa;�D��G|:Ţׄ:������ݿ������^w���!9�8�g�V48���" v��Ndت���/dO�� &�>��b?��(�⪄�㙔�q��@���(�(���R���W����S0�~����@)}1����&�@�T�|�RL+?'��f��ϙ��LM��A�L����V'E���_)�m�]���������a-%a#$�hY&z��S/�':���bj�sq�m��W��<tI�Z��S�ުdT���'���q�$Y�ؽ]�_/�3 A�s%�?�w��(T
)߉kE�	Q"Q*��ڄb�s��(�w���p�BIqQ#���0T��F|pG�t��� �d�����y(_&�u�;ƻE��EƠ������x�м�\����J�恵=vQ�����9����N�y�U!�aM�^)":��w�0���%�Ǧ��a�#z�oPւ���I�}�8u`b��Z�^�ڒ�g+\WN��u�/����Z�i���µe�2�P����M��=�ժ�R����u۷�����w?9>#�ΒL��#+��]�&�0U��jCP�wP�g��p���`�]s��IU�8����G��0����0tTl�����������U������0��HR�2�H;↩�z�v�6j@���ڿȽ��xs)�n� \���cl����94�hqGk_�g��$˥Y��Xv��Ư�{b�H�e���w�e/mh4T{�����z�5��_L+*"J���^ٳlJ�*q�鷋'���p7�v�1��v@2\����\��HH��E ��ޤ��>��P{��r���%�0��|�A�y">�q�K{��D^�w7���/�m��쥣=�(����~Ӧ:4�� A,���R9��6��V�O�q?�|�/��Cz�ntq����9���7�aa�U��b�*dUB��ښ?wd�e�p[9��4V$Ŵ'��\�4Xp����Rg��1({�����bFO:�	@R�}�br��y�d�$��V���/Y歪z)�.�Z{hH��tQ/��w[ʪ(2SU�s�5�-#vG����\��X
iX�uCt�[p|5��
�t��D� �PL#h铣�d�ɯ%����2R1g�����ߞ�
"���W����Ijdn�d����&�C!4�31G	ّǮ��?��~g�$b�m�X"��x��(M�b�r͕�w7�$�r�Ǹ��L�����D��� ā.��ߖ���تeZG�x�F�f&��5��As^�������J�r�$�:ϤI��b^)ga�[�ؽ�����M�lӈ�����iE��_`@�<��K �{e��a�ڐqe��:��Oꧽb�PT�I�G��sN�r��^��(�ຯ�$��L����n�3[�hP��"�&!1��B��l�w+��P-t��y�fe�&N���Vͣzx�Y��#���:d�g�C�\ ��/���p� 48��S��?�L=l���*��vU եfg֟�̃��U~���h��xf�K�^s����j�"������9&�x��Dc� {���R T������w{hW-�g���!%_e<�k�^�`Ϋp��Y��7�ѳS��F�r��J��0���M�:�/l����C�� �xv��5���p	���^VъMƱ�E<�.M�0"�����+�f��*�*]I�AS�E'
�ʺ�Y�����2��Y���V�9��9��גt&{�gY+KKSe�i`� �,�n[�.�E;�֝������������~��aÄ́Y#Pcsz��bȞ������l}!j/��-W�����e���.A���X͜ �4��5��$d��囖�ͼ7ܾ��p�>�9�x���X���nd��k�W�Y\��f�����_J�9OE�y�
���\u�	E���뿘�>�Y5\������o�fI�1��2j�Yۋ��o�����T/&�\��F,���3�J:�JsN��6 R)�x��0��7���LHj�ޤӲ<r3F ��kY'�� m�����?��4��)H	�s���I\�N�I1�YLXBƬ�C�r�8@���	R5�A,��--w�g�{��IB�n�*�eEb�|��0���~ڃ+���e��![��ӌb�r�z�A�=�O���|��ѶqIj'�����,d}���-�[;P{�k����f�hz� Z����Ċ�Gc=��p�R��M�t����-̼&�3[3��D�?=�
�wOj�U'�
y>��?��[a�0���,3��/(h��3��о����6~?>l�U�vlO�>��{ł����ޒ�$7��R��F�H���\��K��e��G=2�ajݾ4��l Q[�NO�jj��ad]���!�e>c��KJ*�[�2a�Y���' �6�9VI�Zk�|Vë�Rj)3�ۨ繗V�������=P5��'�������{��&��ӊ�	�`���t�4�||�w��7u�����?��1�#�|2����"�S��.l�{t&�#�7�$����#�ِD��2�f��	mi����ʈ�,��ɶ2��L�&�M��� H��zz�<.t�������؜���h+ml)UT�}R\V,Ci�ق�й��l�у��$(�m��Q8�D��iўKĥ��	Toߊ����9?`�iEg=�O�`� ��%r*]���H���ĚFh۞���s������@� #^�рճ��@1�U*&��l����P63(��D��bpq��V�z��F��϶i�w7B������.�<\>�s�/e�^�]�Ά!��M��b��ڈ�/>|n�E�1�`���ƛCE�y*�]��E#�@O�.�F��/N������%.͓��8r)�����җ��!V$E�w�l���k��Ӆd���b�.An�p�4 �0�Ć��g?�#�a�׸�۠w?�ߩ����)��u�wA�J�j^F<��T���o�Ũ�o �d�o鐁[Z�׶ `��W־HQ�8�`U�G�L��/���1�x���K���J�d��{����V|�j��kL��b,;G\\1}f F����L��L�1����'F?�u��7�<�)/]!Q�}UB:�=�?:�U,��!TD��&D��*���iK��?��v9찙��aF8��yf�K���a}��:�����w�_������� �쮤=;X1G��h����ڬީ�en�O��>���o�M2���-��ۺ;{�7GC�\����{��$��ľ�(-D��;l9�� h�b����[)��s!�]0�����[����� I���U��TX�l�%f�sݜB"�I�F#6���SMv|IVn�{u^㎎��:����M�������bU���ԹQa��B"��쒭f��$��)m�x�H_՝��vD�!�f��+��:[B���Z�W������������پ�z�����-�`�ڶ�e{���p�#ú���f:��+��(]>H�L�]�Wdo���iF&i��ۄ��E?Dfë39�} /�i�R��E�9f�s�1}�1���m��+��p��|.�
�43g�M�oi�\������a+��4g��y1�t*�^V�Ⱥw�k��X<7͂[�ߑ�GLWE�!����rJt^�>�,J�Ӄ���D��о[��J{����C�=w�K9H<��T����:!�Q��$�r����P�^Ī��<�Y�Pg2绺�Hq,�v�B���i�9�^�m��:�:{6t9!>���u��m�]S��N��h�ޚ�ZWQ�ЁҸ���Ql�(����״�F��a��=.�[!��'Ud�j]��ܰͨع8��	qS{�r��ĪFԧES#�\��O�ЕF_���F)*��#s�o��h�������bU*e�j#9��O;ޖ���l��H��t�-����Xt��Bw�z�K��W��}�3TĢ�kHFc�/R���f-��3S	X��b�����6�Y�7A��E�r�i]Q�EWK�+$4~D}b�p���u��X�ߜ �rG1%ƅ�&C��*��U��JJ����s}���3��I2p�0f���:,��qH�!����&��}ݭ]Q~�C2`u8��Ez!dh���l�Z���8�h�7.�:[�"M08�����O£�3q�2E��ͼ�sK,q�����\�ų����ֳ"���p����U���Dֵ����,I��P�d�~��id�ʣG�}�Eh�������Y�w�$kЗ�~8��|�#��j�Z|BY,�0�!ƴ�qn����`fE[��ߪCn��U>$�]W�k���'������!�j�]1�4Tl�_�vR�?C���Ip2��Yuk�ز���s��$����]{g���1f
����V�X�!7v�;��rǮc;��d��r�U��c�/�
Z�����jS'��B���܏K��f��$��,qi�_�I9��޸	q$-��� G�I�� 8�\�PA�]�,�}�}������M���1��mt�j�}��p�[���pP��'9�=�mF��pM> &��:��T���|"�c��^��T��./6���k�PN�!6{zO�� n	`\�����&�L�b��4��Us�T
<��8�k{M�
�8��5��hb��#����{���l���El�B����7��0h�4[c��e�+����D�*����M@��M͐���A�H�yI�J��Q��L��:�Up+>�er�[��qǓp��%����J�yҽ�-�||l.c�j_4�auU�^��}����ϋ��3�b�� �h\��=t��+!8�Ž��3a-Е-+P T�C"_��͎I�I�����͙	Q���� �pw,3��1�i>J s��zO���R�oK<��͋o�t&'f58�nv�H�:t��F�a�}�~��K�b��ޱ���P�n_��1rʝ��®Q���!7�X6�1P�w�5�G�����C>Ձ�O�,$6��n>�[�N��$[4��ĹI��}w�L*���]�D�+,~�iW=$�<�_�پ}�������U=�g\
�A-R}K
�[��\��	�@[V�`�6$2ǯz�H��Ł��� ���������yG*b��	>��MWis���V�ȷ.S[��5v�vA�p�]�8)S}�� ��zIɪڧ�fs��#<�����3����/F�����h��F�TE�� ���p9G�
y߳z;Durf���Ηb�tq���Eq�xR��?i1�/�����K�d�^�8�Y�K�7��/��{�9�*����kO�ZQt�����?7J��.��T��ĻQ�*�t��9/���Ic�h7 	���H�x�A^��ueP��:ػ��t
����|Yɘ{	]+?�X�Q���6��l���r.��������O��[���=L�bi��X
��r_dtD�-��[�F�������6se��XД����Q��f�9�gX|vU����wP�)��3�J���B�O�쨺� ���
��0�0��g����B��	C�:F�e�F
K��N�I)�X=�b�߱�jS��Z�ؿ�i'�λC2��o��;U��)��s]�.�Q���E1=����v(V[���O�Ҽ��T���^���=�=c�O1�\!�I�%�29VƜf:a"&�"��P��)��R���d h?�Rb3ba0��
d�zEp��'���a����`�7�ku6��3j�(�ɩ��ߎn�oY4v���U�A��SrF���f��ND��1�DYc^Lb;"��&������ʶd_�Jf��m��*N۰�2?��<3�:��,�u+�	�����]��,~I�_څҿ��W��X�9�ew#�N����/�����.��$�H�R�rP}[B�k�U����2B���';�r�v��U���22(B8����ꩱN�޳dR���]��L7B�aaP��o±�[__>�+���ۺ{_^�.��%�Xf�"�p
�^4��;$���d?X�<*�Q"d<�����W\��=K� Cfg)��Pk���kl¦��e�}6�VJfUv�7��g&s[[7Z$� =t?������+�N]��|�k'&3������`��ݖ�e��}i�K��z�'�Kۆ8���7k�X��Ɯ��<�(�Mn��D<���l'!�]��5�#){P�6ڙ�Nf)/���Ȼ��vIpPٙղ�!�	�0��]�'��h����U�=m��� ��+P��*څ�)�'�<�7��/;�qG ��f�o�)V��9��4�Q-�r�g �h:�jߺ1O���i�������2-�υ~UeWDHH�FE3g����y���X����S��Nڎ�#�+#���:�@8�Af��s��\��9�l�����?��BJ]�����K�8��)X�Z��l��������6�8�P�HewO;-�h�*�\߿Qe����_n��&��ur	v��L
|�>�.�sȲ����of�NLTl&e��I��~×B{�Q@O{�Pyg�/S8��v��Rs�j��5�����0�l9vo���k�a3=��4�vt$�,d�ܔ�d�18Z�T�����f�r���������i���L�*f^&�����d.��o����g�3�4O��K��.��veL�S��E���� �Nʨ-����5(Kk��q/�(/A�������oa����*qW�U��G��,�����|U8����A���� �q��Z��QyQ.�c2��>�!�Bs�!�4�����XdO|p���i��
�J4�xc(ܩ��f�=�_�"Dkd�젽v��	n�������<�H��E�����|��˛>�3*5g��~OڏTc�7 ��k���� X��/���i�$,ȮW�:�����'���q��DGI��p�/��ϒAP����#���y�lޜG��@�.���@�l,숚�t���"ێ�x$���K+v|r��lz.��$*��f!���j�6�
7S@9��;l���K�O��}��'B#��kU�-�G]�B��"G�΃��~l-6T����-k�(2�)=���@֜�[����B���X�*����{%������@(��ؔʾC�F[�]�EG2��dM(xxn�����#59�+3 �~�b�b��p�'���F�;���#����E.���M��M)>t����CH��.�����c�J�Yr�I����4^�U��j��AӽlUvn�yS|����=���L?��Q�F+-�_��O��=ת)ُe��;�=S0�hr�� ���g�-ӫZ�,��n�L۩b)��g����e�u��LzAY��j�6'��BRƌ#X�D�l��z�<�o�ј��yh�Э�J���O-�	8n���@/�q�����C��GY��k�4±<��x1��!����Ì�h~��P�t��]�S��WOgv����#�����gn���d�]�g;����G�dų�"��Xf�����'��h���;Tg�T��C�#���D�Wz����Ee���R	�d�Wp�l�P �N̱�����s�{��d��1(-Ԝky��9�l���}B\��Be��b1�V��4Qh��Bw_Lm�c̓�0���׵�^��?�	� W�e=*�@�9�X,2i���Kdbpә�"2ɥ�+}n��t�#��޶�z&A�bK���X�j��[���V˸A'�K��=�98H0�:�T���;�_ȥ<�X3)e�=؉Y]�U��c�RO�	�� gHvV�NO,� \5��[�JY�ެ���Zb���ħ�m<p��B�v���E�|ךcK,����� �\�AM4����ز�h�������tu۾?���^0R�̈́C�b��$�se���҅�/��CZ�Xd@�q#��@��s��+\�}$��Z�o91I�i���G�����e����V~����`_�;c,LCi�#p �]=���4�5�#)j"��p5N�f|?�ԫ!N�)���`��>5n6�w@����ɂc:�n��:EBJ6��1Ziԯĭ8@Np	
8P�����7��:�������2^�{m�6�Zb(6bH7x�udZ�Pf�d���5�ص���&w8��d���8ք��C�>��|��J�?S3���h;��}>\�@�z�qo��fz�����2�ewR�&�^<�5���7)D��u�w2�w��a(�G�fo�i��B������k�a*�@��GF�q4ĥw\�h[nh�6F�n O�2� K������haj���Y��lqN������PC���v�F��e�<Ƨ�d|�/L��͝*K�Q�t�~[�x���@M懚���	ᾜ���Y���)�B1�^k﬚:I���[ *僅�9���!�+����7d��X��+�'|��]u��(�&�9}�c���\�H�.�o�<��>n��g�2Cuo��F̘ix�GL��פֿq�:P����]����(m��M���{/1�#Z�-%�\��g�{�t_43 �)�E��T�����z��*֑����.�/ظـ&��I��L���I��h�P`P����k#������Ӫ�$ B5�<��r��
��}r���^��ᵯ,��v�D`V�UR����VH�̖$;�W����"D�)��U ��D���_q]���/�[�Δ1}�V�$�e��a�(�&����U+5��lO�"h�����¢�>���D�T��0i\�l- �)$�Q>ಞ�:���|/Ȭ$��Zi%��"�c���3�^~�\�n5����O�d�����dDp��N��۾���8��f��
o�)]�(�.|�#�
��YVJp���7/��!�]��!d�������i�q�����_ A<��ڽ�'�<�N���Ѻ˺e�(G�7��X��e- ?�d8D'm"'�;��ƶ
u�
�u�yM_�3����J]��*'غ�xDF�މ���Fۢ46��#ԂX0-5*68��	j/Ҿhx�7|�g�5�8zZu/�ggwg��<譑��i�Nx58m�?���V��?,�v"N�i���oZ�����':d��kw�=Dع*�7�w{�|_
"v߳�~��]�f��V��V��M4�Mq�.���_Lj�Z��U	JTW�pջ�����e����tΑ�5r��n����y2�x�o#�JY��4�8F��F��W�dY�\�#���JM�W`G܁]O�D��WX�����t�j�?#~����a�=+�O����|YG�
��;���Oq��v������g��LΚ�>� 'O��K���n�8g.��l�J�ا��6������d�4<��Q��Sq�U &��
�`��g��qJ�E��`V��_:�nH���)�0�te
2��.���
���UKAĲ\4������瞩KIʁ�@坎'>_=�K#�>'K��+\�$ϴݠ�~��m�#� �J���:��gѠ<�1X7o|���N�Mx����>�pT��9[T�\zhe�,�F3�ﴹc*|��|ZJB^S͗���ń���DuL<��Y�̈́�Ƕ��1<��[O@�I`I��m`�H��V�����&Ή-?��P������R�Z	�S��etY76�oa2�-/�[R|�{�t'�6�j��'�B<X)K�k�y]�n�������RU�>�V�=����E;�iol�P���� �;9k���|f�z�7M�]���l8ɠu�s���E|��R|?�4�Ҫ��J�c�'�|,d�}�ˮ^ ���C�Aeu��[N>(Wb�\�:���R��-fu� �M�W����6�ԆI(�W���4*��Y�(!����J�و:�����^t����8$�u��?͓F[�g4��^B���[��Af2j������_в���^m?<1.����%}�Y�8�5����Dmuw��&&թˋm���&3)�5ұ�`Ѳ��Eo_ߛ�
I�D�T�4�����)$�S��J�؋NM�Lv<1z%~�$�T�e����<� g�Os[?��]���ԖpI������:��m�~�_"�����{�g�Cjё��;����I��3�۪z�}�*��4�"�0{�O�~Q'�vl
��o�!4T�9�1S��_l+��T�I�k�Y�i�ek��\)�Y;����Bk��$7�#Z��H�D�pOW������޲��O\8�QG�/�j���i�भ=�� X�̔��h1�BDD��y�p���-̺1�X<_��Rzf�ݒ(M��D���yh����<=D��r��?iD�7�
X����0���<P�m�-J��Go@�Ʈ'��[ɥ)G��m��ڷ�$��Q�ɖF��O�,Ƃa!:C��I7vaQ-��Q��&�5d��o����0�H&���µV[u`�;����bBu�҂�=//�5 F3"d��5[����F����u��s~�o� �C�FI�9v��*�֛u��_r �<�5�����r�,a"�.�!X�BQ�I� X��9t (TV�MM�@X�0�oN��8������HRp{��])B��ݼ�o1��П�*LD��e�z��ꉮ.O!}*淦�=ˬ~���$�����컒�D���mm�\���zf�ԗi���]ã�����n�㠼�g)w��٥:k�ޞ�z�_/fm�j��Ќfzx�ʈ�����Cī�v�1���`Թ��e��*}�]�'p)��S$qc�j�2ʶ�ך�T��:*i���&��z�Y{���g�^��-��F��(�H���\� 0m6���є�(f���qC2|�M�.D��T� L�[3�cٜ9�����Xޒb/3bQ�G���@zz��V���C����`�78����Y-%�`o�����(�lh�LVҞ �[Lβ�˚6�L/^`J�Z�QYV���gA�z�
�*t���OQ�lsaan�X�rG
܈ho�J�⼣�@5��^�&��s�j��"W�)����a�C���g��p���Ӵ]��y�ʰ�K� �@�$�7���%Bp�^��w`�0���09�7�Ֆ�����{0w�����?j~#B;d�K�Y&8夙1�t�����% �2�$�?��(�c͆'��ҵ�q���;�zi��/CgUNSq"���,^+w:(m@e0�{��������,7j��O�D"R�e4��Ti������J�r�S����v+�򏶙Պ�!��s��fuY��������p�Bй�/�3�f�s�.]�12��w��_����W����H�E�o��	�׿r�;C~��%6�"W�{�Ę�)�[���󉛨x{�7~W�H�t��\QWÀV/Ġ�t�v5C>[�R�ⴗD۔q%UtJR��	H��c5��I��=�j�N��Y�we���*�@��O�3"��4<ޜJ�u�m=uj�lחu 
G��ǲ�Nn�XGԫ9�$���7��Cf��Yr��܅3�q�:o���I��ѲR��o���x��!�1/F��ٜ$(B[?�Mf���U}Fܻنi���&�+G��N9�����ф�6�$��8}96��s�M)�S �¼�cN���@��g����n�/H�H{Z�v����>C�}�@�Y�o�����I���erW}�#���oUƝ�ߨE��:�L0�#I�xd�h����&���@-ցƖ�A��~tY��<���1C ���ub�0�l`C�_�ݣ��HGQD�9���~���	]�Ӓ	�.w{; �Z4�ʓ���Z����y/Ǧ�:� \�1P�~{��˾"wt.�FS�`�H^�0�f&��nDŁ���'�@nyc�"��?eg�U�Ћ�7Z�d�~�ޮ�Vio������]]S��R |����K��J�}�F� �eW�%DFz�)?X��F�:�Kϸ�x�]��N<�X��jH��vN]_���4∯�zx���߾|���+Ǡ&�W?1 �W�Z_TN�v���߇r�njxC�b"�������w.�{��e0�N2�z4�w����i����O�}$?�ĻĆ���{�|�t����w�~� ��r	CǶI1�E�A��^}# �I��>����Ő�N��Ӑ2�QA�!���{�Pd{&(j��l�"��Na{����'�|z9+���h���i��n
�_�5� ���v���w�_��	<� )8r�,��P2S�88::v��0*���lm��4���s	k﫣.lS��zy�4���	�c�Q�&jM�a�6��\�Ls	l���f�������̢�n�ޏ��;v����x'�����(e�mt͸�>�'�-�[w"7��;��D��4�I9 �2�1�#3���s$�ǈ�`�