��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�djB�D����)E霐CJ���@���/�6��	77ZP �y�0֥�U>n���e��� S���x9��`4�������E�ynT�t�r�/|���)����ы����tW=�������C%��=�1��B7�۶�b#�3��#'���֒5b�v7�n��)iiWw�a�~�	�]�ƿ�hC�KB��L�mͯ'Jl5���'t�ss���o8ױcL���j���4���i����������>�OǮ�	+ٰ���:�h�3��)�tϡd����l��sG1�k#��S�K�qG,��+����RĲJ?G�G��n��U)!α��<S�/ٯ�*�����lT+|`���ܺS7i������\<$��8��2>�Q�m2]h�Q�\, Ȗ[$� q)@�UCNM�  ֬C����?�?�hn�t�'���	4���%��z���������'�-��S����v�9�s4�z�����G�?�f܀C�8��0�9c���kl��[^t��a%i�=��0��'�-�/���_����Ոp�F}���ۏ(n#�X��7�0��׀z4����~���	�cA�r��@̊r���ܤ?�ىM���DyPR?�/���K�}����^� (�Cf�D�܇M�k5�H�(�p��M���f�k(!Ҳ���1�~�jh �@��	�H�,L��B(��%6V�u�niS)����[�;�yTc�����	�n��6���������q����H%餞�����M��W�e��"��L����P�&7 ��A;r�}E����)���<���מ���mn=yFA5&��ضU7_RT�V��\~c�OE5����u+@q��T�c &�,r��ˊG*"e� ���z�7���X���S��
��tC�3$�2g���D1��[�;l�`�F.����[EH�m?����ں;䠱%A]�����v$V�;:#N,+{|��(r��<����U�����ڻ��JNЙ?*���|�*�
���{Z2��x�0�eDG��u�>��:���h$��,�:Ww�L�^�7�'O�6Z��_#�J���܆"EH=�u�d�ct؜���SS��r��a%�*K�b_Ι�����j�gW�cD��U���%G�oF�ôx�|�(cf����j1�� Ur���x�,6�c۷�z͡\��
��T�zN{ش�N4�&�8��e��c��[tl���Z��F�����zqC����F�)��U�/�]���0�1�2����@�!#��:��)s~16l���,���KFq@�t&���CH-0�P<A���컬N!O�����I`����_���٪f���͉�E�܊��=I���콷������ߵ�+�y��ԣ�n�
ְSօ�_K�ц�V����ْaD��>��/lԾJb�~��^���'�䆰��,�����R�j�Q��it��/6�R/<fRi"ބzdw�����^6���g�4�;<ʁ9�m)$΃�#O(q�cR��PT��3���m-����p��?��0BU,p��Y�ws�J��-��ͧWh�a%�����& ֒��9 �ϊ��蜔*��rb�b��0WJ�mc��ڳ5nz3�W8��G1�l�������h�/��1��K8���q&��.�R[b�|]�̐�x��%1�� �ĩ!9�l(@|�+�����1IƏ
�R#G����w3N���L���?���w޶�f��	���KG��U�*~�il���
|��\�5�ʛ? �_:ѭ|�� 
R\5�7}������]#&ז����a�56��Mj�áS� �7]$��S��b;�\`�S���s��wc'�ʜ�����<e��U�J:\X�����ɲ�B��߻I[1{5���'�����@�`�"�a�K@�-�>�Hw˧H��r�$j�п���k�\S\���F���fI�EM��\�|�85D�B��DN}C���X���Sɷ���lȦ�!hx�y�j�O`6);�,j�"IB����d�eܕ(�0�w~�wWĭ�;_.���OH����UB#sH
m�շD���)h�����%��oZ�ŠYYOԚDM7�Жʇ��0+E,�����`����D��,I�vܾ�@�K�ak��t�͠TI����.���ͽ�}�P��K�L��Q�.>��P ״mX���I��V���&R�8��x�X�̞�5��>�$��eBy�������BҦ�,"$�R��J���y�nۤ%���u�܅�{��A�Ĺ���q�qk�	��ҺG�;��L���<E�7���BVrlv%kFl�.�!��߃���r�V�O8`���0G������Y
Z�.
��rWk�j�t�}p~=��Ǡ�upC�|Z�=�W$!k�2��'՗��L�%8���P1`��H�4�c��d�x�g�Z^���H^jw-�t���Z�w��Y�H-�A���zh�o9L����G�֡�.��GC߉�U�i1��=lb�/���b�L� 2B�\?#�8
����������� ��@o�<N�ż3��k�V���C�'* 2f�ǵ/�%M�lg��却���XN�U{�gX����2|�y[��Еj,�+��`�'2d_aT�D�ƪ�e��(���dƝH�H`�ƹ���V���T�~�S��Cаt�#��TN�w?$9���s�+���g̢�ah�z�f~�
���@U�6��'i)���׏�:`5^��.�F,>�:�eE�#��?�X��P�SEY�!�N�>��
m�M.?��CB ��L_����DWr���p:?%\cZ.�ⲙF}o&�&#����,�֡��^��m���V�K>qH����ț-�.��o�z�9�$�g?�^�zT�0bS^w�
����/�.��
6���8��-�Z�W/���B�0�:x���zM�I�1�+�ݱ3�#�%+x�"I�=�f�GF��6|m�
�
9�,Q4>��c΋ � B_�xQ�RF�Zf�k�������l�ናf|��--ܒ�Vr݅}j�g2xG�q��D{�nF�� }���aﲙ �#�z3	�$���+��C�7�ѩ��/�*�w(<-�A���b��[U����hsi�Ė�W��ŽG2Ƙ�4{�n�#7�W�`��S�D��Yr�.���w��;��~7k���%�g�bSsavY�-�-\�.P �p�3��|s)tQ�7�$x����f�>X5����"������h!xG���G�:�D���QBtOc�'�ŏ"v�\��2�ߵ�+5�<Y�gi���v����{G۞.+�Cr���d&5߇2��ےE�%�nx#/?�Bm�����ʚ^u�8��y�<��r�_ѣ.*r^4���aPjP��*ChB̷K(�'֮ƾU0őN/}ԕ�jn��\[��-����6JA�i鿺�2h�"���ᔐ Q��� �+p�(��S�hQ/���yu�ƥ�]��]��[�������B_��(�Ro?�hL����ٶ��,	��s�
�ƖT�F��O�N8}b���yYӫ]SR��}yv<ۥK%��48^�Ź;��%,�Zs��5��޲$+ێ�|��7E��)y��Nw�� ���tf�t2�+M+��g�f�����n�����	���!W�4��eIf
K�xsĐ5�$H�QI���em���JO�坠?`W���_%���5�U��+�(�x�?�C˜�lL�E�#�.8�z�̏�s��a��ďY���A}�֊�����-����w#L�G��Beo�v��N}��o���K�:�>�$�SY7~�	4GVz�	����EiZc�)��g��`�)$���FoM�X<�4�H����^r���7��y��3Y,'��v
d��7���'�QV�s���Y����/�X�a�.����伶���ф�p��+X�tb7�
��o!6��2��>�P�QA��q��k^�+����
N��؆��X�������G;fa&%�k,��9�`�n�Ma��N���éܱ��7�I�c�BK�ua��8��L�hPF����ԯ���:ؽ�/���L���`�T��ݲ�𞩆�G��
���s����u(`�������Q��O`Fd�TNKBi�