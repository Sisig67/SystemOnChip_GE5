��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��.y8el���SN}_e�*�x+�:x�@.��{(L���i>�*�Y���f�0tCP��l8H� ��&�l����\��7"-�.kC�ϕM!��H�O#O!���hjf���5k�|ENR1%��9�R�"��5��z�uЁ��2u��9#02�W��=�h���]�n��ǰ�j4����u���A[��D]���׹��AaMӦG�5�
�x>ʭ�CF�;ڃb)��������];�<��5�I5^�mFO��𩃈��c���j�X�Y��œ�*N��N�|_{�����3�� ��#�O����������6��RKJ����w�ȣ_(l�Ÿ0cl+L�n���r���}�m�'�ug��K3�;��ު(���+6������!*Xt�y��j������@S���)5�����B����`:���d�E���wdrx�ן��U��f܃�N���_��3�-��΃g�^���X��S��R�"�q�G�������t��֖#g��݋�^����!5r��v��D��L���뻛��)c�wp��D;�������"��aadߥ&A��8EB���zVg����K\�!�:pb&ֿs;�ޠKr��YK�qf�f�.�g�n��eК�"�?���ӹ��aH�_���U�|��GAݓ���$v��'��'b�.R��7�<�2����v;Nֳ����?Gu�݃ęP6���"�>�%N-��N���B�3g;嶠s�!�m����
��E����2��k9O�L�͠�h�Lƺ�pj.�����S��� $|�n���Th�*5�����ϐF����;M��r�qb�<Ǯ��8k��7��1"��B@�m8����
���گ��؟���t�Q{��CoW�e�Jmׇ�,5�cT��"$�r�:�`�K?��2��5�iO��RN��e�Ƌ����J�>Og��.��(�u��@������M�؟�.\MdG[U9r����Jh����-7�����Ck<3Z%�Ġ�ޏ�(Z�)>R��'�4�`���������Ϝ���T,��t�V&K\�� ��G�}��}��)�t��8�Z��>I����Z�����e�;Q.hϿ��/g�$@Z����^�0�E���z�����Ic�:���;�)Tf��EA�o�2��C���-�VH��G���%㳩�L���쥝(�!ӗ
��&�טu˥��4�ݘҗ���Y<���G��w@�����f=��Cr���>���LXp;��v�L��oc�7�����O�RQHwc=<$My&8�����n+�arM,�y/��.d��8���X���kT9xfbą�W��Q���%�zI���z��9 �4���鰑�զ* )`�e(W}�m�E�[���v�O�<sTd86�nW��S➸��mO���Ҙ��I��	��Tm����\�{�@ča�f<��O�GY��_���=�|�8�}A���!`/�K�E��_J�2��zH�V��S���E�z�P�	�`2���-OĠ,Ne�&݌A��@����Y^l�|��͏8��v� ��)���5���GO-�~��V�Q.�$��b��z�^���v�jc� �c���O� �$��0��5Lmz��>�=U���?�#¹Თ�[�ziyfC�:j ���|q3�QQU�b��PA|-M#�h�Z^�M_����L�w�|!��.��m�x&�XC1&�T���}΋_N��bz���8ê���D�TJ0BE'1cu��������Qc�A �����_͏X��X�j�|�5���9�z%~.)m���Φ7��	����=#Fgz��rh�Н*F�&u�Y�t���|)�"��]IR���7T�d|��r��5x;�\��8�P��<�4�����)HdP��r�pJ�J<^�l|��,r�O��6;�IS�@Eud" ^�z]F_�kҨ��P��<�v�v㎭!&���F�j�{�šAv�O� ��d��e�������uT��ʎQ��J���ݦ�k���Ǝ�X����TEd���w����-���-��s���N�8�k��t��YD�6DS9��_�^�
 ��.��:+��?FX��^�m�x�d�1�.~��_2s�|qz׻_&t�3��KH���R���Y���j�^`L�	ʪ�[��K����XG�7���c^:��Bx_Ig1T_�>Ѣ�%`����<��_e�����*��c����&:*��1�.j�sȆm�Z.�hH��X��_ܠ�2l�	@J���l���Li�[Y�W�솳� C�*�D���.�0��8՛û��p�_��  |��w�O<�}~­hRW*�Yҥ�Z+}�L4��*�7Otc�(4���Zl#��ml�����6��}෗<�C7I��m/�E6�Y	��S���<)�^G�E�Õ��}�{�����q�@���0���+�K��¦��v�pL]��H�5K߸	+�v?/G��Nc��Sd3l�K��κ���T�PU�x�-S��4��_�a*�Q����;���d?�Z*�l��[����|���