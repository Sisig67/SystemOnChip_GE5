��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���!<So���2��E�!�7���feI�R�34�F�\1uR�XO.P㤳��"����(W�����Y�us�'�V6g{���/�Y�^( ���Ne�[�����8�1��{SZ�k�eZɇ�FUHn�i!�kO����r�o�40e�@�̺Na|�g|�O̲s����_�oW�h+c�	��x�1C5�]�`��P�#�Ι��;<��C������^c�4�\us	���S���x�~T-���]D�lK�c/[G(+ف���j�H�3!`��|�V�k�)j���Rrj������+!�m�iS�\�,�D nP>�:V0�(�9��O�Y����m���7Ӧ�J�Ā7��-�o�6���d��iP�2I��5����^��1֐쬳پLƑB?�(�x����wj�j[p��ب�Q��8�)���b' �{b����Z�مIt<8�3�\;++�Ҭ���7���$5�?��Hf���*"��6u�Ea1�Q�g=�f	����%'(�l6���g�L�YG9�:x}�� ?d,2+5���1;T��U��Kڐ՛vN��~ō능���d�>��$�s�D�Kb��{��V�L����+��6pM�ld���v�0f3���w�ہ�V����W��� TB�Ov�4T��9k�m����Ҟ[Cṕ�Q,:/I�ff7M�d�$#*�=չ/Ȋ?@O����-�+�g`��0�E�΢f�Ր�#��l9LBi�-�.�{��޼W��������Jx�a�8T�r���ŲG��@�.�f!`¾F��^~�G|�v �FLN�j#!Mʤi��ɘ��R�������L�"��[�V:�(V�R�Н7�i&O��Q3��������>ac-k�cq�"B3Вa���-D��+�;�IYd�xޱ�T��F�A��Ji	���π�[�>pE�����ðh7�A�P5�f7������:��_m��\󔊁��?<���5|���b�P$1u� �,�U�����Q�	$��/s�QC��Tb�����nO���n�E.�|�@��}�"�^_"~B��F͵�U
�Zյ'��^L18ik?p�:�yo�K���&Q�V��b�՞�	�Ja�2��ň3�����c�R����k���+�T���0���A�]��7	�*w7������2y��� ��#p6�ݴ�7̧��[CEwEW���ȴ6��I$��Y�Q�[S�>2D��l�J0�)J^.R�ÈW߂i+t�[�J@��*����bc@�8#ɠ'�gu�5��eN�������2	��ո +�g��bC��T�]�F�l3N|;�W%�� ���S�o�,_�pW�s>��*�. 2<*���s�7�����������SH���8�8��I��L� x�@����`�M�%� �3���R�U�]�%��N���C�x��ק���Yu��3���=w�Q��#�"�\�qʟXe�?T�4!vd�5��Rw'0:��% ��V�����4�X��;G�O$\�R
g�7��D�x��^F���p�����Z�:���/#vz}�xנY>b"	-}�v�s��D�L�MŔ����C��m.���P$��8FL�n��Z�r�FRV�(�����q�6P��J�b�;�����\���D`X\3�@����>+�����ow5Qm^?)]3`�%B��36Hj���C9��M�Y�c�7v���x"7^NJa�\؁��e;j�%��U?�qN�룂s�"tӄ��H0g�,��n��D���DŹSw���[��1Ԇ���|���1�-i+3�u�.k�_L��!�8��@WĚ�)�D�PoX���t��wK3���-w��ՈZ�^�Y`yt���ƕ��FWry�E1�n̞<!,�FU_0����\�`���px�8 <���Q��p?�+D��}__7���'xo�X�+;Fh�yt&Wm;b�}ˍ7�C��햪>��}���G��`oOw�7����8���}6���Ԗ��K�����6�i���I�+Y�~�J!r�5���G�90�~�� t>=��@��2�6� "�C@F6�� Z��Z�2�a`-�x���ZLKp3Ǻ�I�M,$��ڝp���^�zzn����ĺ��}�b|T�E�2w�B�Y��Q\�>�
6~/<ͪ��]���� �����j��1�H�l(��{\O� �Ս�S�"~6I�14�\*��R�ᜣQ�� L���3 i�<��
.���m����sF�V����nT�����j�?���<CH-��'��~��n�j�&�9��o}^%�p�;���4��;�~�(��Z�K��3��~�3\�=֥�l�:&��0zLg�gipC'�s罏��ONj4�s��!'_M��K���d����Њ���B�܍q�,�%��o�@���X_�Z�aE��q����������=�;���9��ǔd-��҇�Jq'�0c8�DG�ut��rP���X:j�#f���4���٦�Ɇ^%5�����,�1�����\".���;x�ZM�"
.��NM�aC���hs���*��Mw\�'{��ʦ3��V�-�V",,�@�G�+Bc��Y�X^Tq�K�A���K�;��9�zX�夥�Gi$!vI�1�2�轷��i.���dT˹��e/\�%�S�E�M�N3Xk.�t��6?���n/�<#x!D$�+���Є>��U�BQx����b?yL��0C��#!*��:�9d!�i���#� {��r7F�o���!��QQK| ��d�68�뜋j�	�~F��,���ʠj\]-qψ�x��~����$*T �pn�Mx����8jyMz�n��:@Mg|<�
JEU�-3��[�q�#�5b��\�h����e��.��<[�c��~�Z��s� I�K��w&����B����V�g����w:S���K�_���71"�Qs�𲰑��3 b�Fr��A�U1�\d�e�����|�Ĵ��}��?Q�*�IUf�3{��=/�dR��4�"ϙ��o`D���(�B��A����n�Ē�(7=n�<�z_�0���^%(�@�@:�*�Q3=��[)&8�1d���6o�}��"b����+��k��ٷ�m�n^�o%��ݰ�������[������'.ZZ�!�o�8;�+�%�xi�&���T�;�@���Zoe�>0�g�ݿ��ƒ�}g=���pX�"�U��҂Z�ԇ��>ik�+*�%+sm�(d��뻝��Jݵ#��U��<���D�MMd��� �D�Q�=�����G�y/IA��/c��e�O��
lL	���8��:��H&g�D
���Ի+V=׶Ⱥ#^e�C�e(gzo�t�������K��G��: ��pTη��d< e�)U�\�"��<�aX����Y��!�(�lG� �������e�>��|��p��q�M��ŗ����
�nt?�(J��2!`=�ɶ����p}o,g��L�{Il�V��_g� ��E�~+��_�z������s�!]3���I�%Ͻ`�j�A�����q�£c*rGq��¤�tS���N�׿���n�0D��Z�_�,�����^a�R��;��e��Hh��C,������� �$�jeL��-��6��īi�Do��v=j\�`��~�d��p�Ie1�%��6�4��=�G�����z�v��P���'�k�s.��>z���O�A�XPطK�?~>	���H��x�uarpmrOе(�C#$��>�KLPʭ��Vs�e���N?�`�>�~>2]����Q^M�z^pd����k�q�8���l�o�R��������S�.�;�8Lf�/�,.��[��4�y����	2��Y\������EC�`;ކ����ؑ��1(����%�3��*x�/jw�`&v���-�����d(�B��p��s"w����,A�&���.O��]�zV��oc�,���GW��M�5f�d�����:���S?��K��P��G���ū�xl1��凄�8�)�󓵡����4p���=��㶦-�d�Q�R�5SS^��*�ަO}d�)}��L^��O*��;��o&���/�Z� �mxh�n�3캥��L��U@kw�|܁�%8�n#��VN��L�d�]�K*�f�b7�U��=|�,4�@p��3B쩕y֚|�ݝ�c�U��y��/�i�9� �>��<Q}w0w���|��L�P3G0#���
k����nW,ha���Xx壄-�WX�=�%S�
��QЯ�u]��Փ��~�FU�Nj���9�"�+Ȳ&%�͖˃~��2Lz�Yx��|��^�3��� ��3��_k'��K1��������֋��3o*\�鰔�ꌦ]8�F���-�OZo��[<��~�����UB���f��#�u&� /i����A ���+;���X6a�����#�Aԗ+fE���I{��\+P�uz!lD��79_U�V��cg�`+��x?�O�qݻQ���	��@�҇�j"��8Y+ ��l���tHC[�8�ߝc�1���Y�~)b�k1s"nG��u�K}�p$v�A���� 	G�$tfI�s��O4[A\����	�.��h)��V�M����[	���Ύ�A�����H��\M/�;AƟ��b��g��Ϻ{�����3[����]�Y�\��A�>�-���:�`��E16�(�r�~���|1u}��:�����ε�(�B��ـ�����	=�[�i�o�d��靗k�y��(ś�7dp�M��2�a��ә��0^��xI��f��ia����֫�����I@uF�d�T�F,�z[+��u��������ք�K��A�.1r�U���QBg��sʿ���S�@P\H�r���2:_��Q����&tś���:�͞X��U
*�_"Wi�=Sc�?�;g�����,�E�,�Gf!��)�;����&>��V��I`q�@z#=a�=�F�4,=j����Pw�J��tG38����m��a��Te�7�-���Q* ��s�3��p<	W&��^�{�PO�\h3b�Θ�%�T���h��)��'��B���-�=�1�oAOE�K`y�^L��בZ�5���i(J��t3���"����t�I�
��}���+��PX ���26�1淠
��A=�d]��G9o�W��:��Ca�4�(%�qo����S=�q_���@���`�b���Y [jl-|G�Z&�Hā��~c�t3����$�V��17H���sN���a��=[�ża+��E��(RȬK����(
����0�BuV�5�U���!�_���@�_�a#v��*�(P�z~k�9�ZH�IR�ւ�����m�V�r��hh>uj:�E%THTPp�� v��6�ӳb�_�$M���k�窿��'�/�HmSci��ԑ]���T���$l���S�B�n1��w�8�#߷�����XH2;�:�9�k��
�Q�z�00�����h�JW�F;�Q���gh��u��ϯe�T��>L�G��<�] ]�Jf�_>Ί�t��aA���)w�����'��L��2e���͍%����k�ү���k\(���Y��N:/���1�؄�h��4ߤ��z�c�[�Qrӻ�t�8�!.�&�՚"��nׅ[-�e����>��[>���yA�:�PSiQ���l�A���v���ϕ߾w���N�m���m���`�Mj\�-ɒr�|}~��40�(m�� K��e8��H����#ԙ��(�/ϔ�����:�K�6�_33�H���S>�A;�ݪ�:?,8.��UH���^z6��t�� ����w
f����ߊn��IG����u�lM��g�̎��`�R�;*}4����r˫��]�]��r@�:헞�㧷p���7hX��c
H����r���%^�[�܄�;�V���ͫ���6������K1���Q���Ծ��c�����Ad�L��<v�6��x�ZD5�㹒`����	�|?��+8�IE�\ԥAu4+�x��������:���*���8��0�/�,:�7�u��G���������C�n��z���/ P5h(�u<3<���w�4#�vZ�����<MѺa�#�����u;:|�i�6�D"��w��X\��q�(�N�&Ap$��>@�����ʞk��KuNp��C�C�JDר��*�
��u	֭��kK�e����i��i4S[W��G�d�y6��)|�� ���T{(۝�6ÿ�sZ2#� k4?V�O,_���sҩ�Wk�n��{��1=�<��`��=���0ju��+�.�����L��`�Qt9�ܱP9;_Z(Fd�lx��]3��-�eCFp�^�����nwH.�_bۅw.�ʜwɁ3]�����]�>]ΖQw�z��~����J��iX�l# E}&F �����ߘ�F��2gsk+{�)��ڱ���?�]��3�R�!0�^i���|Mg����PWl�Z����wt@7�%3-�x��WP(�G�p��I?G���N��1�F�i��V���)Q�}c�S�2�dn~�*�ez���o��g��0�O$� 6������)Lx�:��	/��zHn}��,ӓ���*�=t���|<_n���_ZQ�L�f_O"t�HhH��'Ya3s��<��TE��9�Y�y�]���P��$K 5�83$x�G}��� ����n����w��,!(��tR�,�VM��.�MPw��"�����H
��幟$���^����\Rn�5���C��s/����}  ��oA׽�e�X"޳�BS[��X��/_���j�
v�W�-�+���x�6'=cxo�1�M���잁k�B?��-�O6ݶ�n�����u������n��h�D4,"�f���8��L?���i���1��?͙���ފ�����\䋙OA�F�Ύ�����.��L����d<t���ʱ���Kҙjf�1�~�C ��E����&*�F�٣�>kN
����]��D �u��d��c�g���&�}��5x�3�їk���ct7rnT�wE�����Nv��t��fu쵫#��_1Zq��U�
�}�N��+Z.΀��ō\�>b�'jS6��+��cH�פ
YGȢ����T��j��
�K�&����V<���ɲ�\��%��}B�+9eEI�_#~�Mڦ��F2L�tP����s�K�6���9_�}�S�'�`J�ϛ�Y��t�5� ^e[/��bl\
O8 ����cJ�i���i/�|j#~۵����Y��e����g�޼��B�ޣ�3�7�]�����>c��ڃGI�˻�����^_�*1a3��*�xLJ�*z`]Z�
���<�T���H��E� ��Ka����e)D�z>�
~��ӗ4�9�EL�o�9�X/� ��l�hǠ���%�lA�yb���\I�B���e�K�px�JCk1����Bc�ҧ�6X�H�V1q�FYx��՘}B������#��ߥ�Rf�� �Rv�&H���[y @�z���[ڽ��� a�p��`k�.�˰��F*�p"�2�w��kb�sn!�n@��Fp��wAz���s����05�l�����y>���u�'�}7��������x�2⬄↔A���b5�`Y����1°����*�	��P-B��֠���_8=:������/�aQ��l��(ދk�h�S�Hp�*�����#� s(TU�0���
� �ǰN�̪%x�0�J~�1����#t�v�������%}������;C�i����9�Pa�4��j��0�Bņ����K�-���߫1E卯NV����l�YC[ك���QD�Y�3wj�i>s�J�TiR	�
��.7���'�-��i�A���[4�0s ����PR��(sK��:bM�\?Vy�{�
:i^��1j�l^�����%��S��z���2Ȉ����@֌ o�v��M���`
�F�+��4�����ɟ��ˠ&���}��e?�#_`��;ˀ�`���M��O��V�۶8�iSA}�u��t)^��	�u�!�c�}�+�!�����Ѧ_2_d�'�C���00���<'���
�I�&�e�$.�N��܏�v��n{��綦���nn��x99՜���6$�Q�|eY17�l���6�������k�{z��Z�g�i�A�a>.�Y��>���8}u&(Ov���zH}{�t5r|z�r������Ls$�[,I8�^�e��I��ӰT��¡�<�/Zo�5^k �Kٍ�����<t�?j�]۞g��M�0ZNvѽ�����%��4v�ҕ?m��3��1:FƩW�O�;J�(�Ⱦ��>�ܠ�|��rd����"8��5h¶�](�P�%h�$Dud�n��f$oe�����i�q�ɫ��>7���������B���V�N�|� ��ӻ��uX6����G���]�c�G�b�I�%ܫ���+5;�-5�o�7���52ZE_��&�Xҧ��\��f�ۄ�Sn�������ڛQ��^���K���鳯���1zo���p)S�V�	e�m[r���Ƀx���$�o�CRr����ڒK�!��6`0����#�[�"�GRuI)�5�k�qZO�\���1<{��[I����NZ!�:���w���x��~���8�f��Ы����v�Ă�I���-�i��=BJ�%Jg���g�ڸ�_�����W%��ޚs�G2Q�����G
_��A(L���'7��ی���z'[���T���#������ 3fe�4�@㒺� ���t�����2ك���O���^�Mq�+���)=��l��k��Ks�g��Ev���/���y��f'@���z�|�Ye?M�։�U,1�b�P8f�h�U�bgd< !����Z� ��P{�6AK���Ց����]���t'�)�a%�R���L�v`�6JF֚�s�E��$j�(JZ>u�p��L�̄�J�'洴���hm�B��['��f3����À^A����*n��F�H=��},��d�L�����\��X����V�w�%�R��8��ڏ'-��7�5k��P�:0����s�VN8-���;��f �G8���W���Xt/Bx9*B����}�O�4�����nAY�O��se�/�s{��n�g��Mw���9""^ܗ�؇��E�"�p�.�;K��.���;��Ʉrۆ>wV8.�E�G��TP?�kzT^M��Հ"�;�$p��,��k?`3������l���#�I���t�&8��	y jehz���S��
�NR��(�XoD�6iZ�����J/4�泤� ��֩r\bY��}Q�o�&�x,v��酪��]vF���՚�\ �N{sw����m8��XP�¿?���T���)�=̲m����0�!��/'T��	�n���ݪM�Aj�K�JC�O����
iw]�h����HQ߯޺i�,����v̉�P���!S�]Y�<�������ڬ��5v�%�/ �$w6���v�'���ni+��H�,�<*���N@�� ϟI�'S�P�~!�%�we{$W����U��d�g�o�M���c�F�g#K� �Ԁ�㩎��Br�m��b������ ��7�O��CM:��� �(e1V�o���T_A�����}�bt_<�6gT�
/�O%x|����&���  �����C[eěm�}&��l2�M3�H�*�q$�6���`���%�|����1���< &j�)����f��6�#�EQ�L��y���gK<=���&{��d� �����91�)8����F��gkgC�����x4��j̊���!PKҦ�W::[�y�qǢ�}�w�u�Z��8�
�oya~��N���2��ݩ~�u{����w
>&b�T���h�(��a��� d"��Ǝ�jT�C�T�C�6j%��뢼�7�A���P+(m$<|=0���
ԟ����3^MK����O����g�fqw��L>�}��\@��n��=4�B5of'����F�}uŉ�s�ׯd�"�	�|�xg��oOt���|�3.�E`T��^�:I`���\�V׫ j��F�3�pȍ��8N�/��:_�IYlk�NC�)A'�p��Bx#�>ZPq��I]�q�:�w��XV"�/X(�E�tMU��������p�v���E�e�h&���z'���V���Bv�Hd��VyX�ؤ�}�S�C��d	�G|��(��ï��KH(Oy�uY̶5�#?2���o�{�*�,_Q&-���w8��@������`Һ ����H�(��+���q��q程�ك2��"#�q	��T���d�,���q,�|����u��j3��j�`={��V���i.S������_䕆����L��I~�� ;�[�Ԩ��5�SX��)�BA�ڂ���MWw�ڬ�j�ɚ�ֈ+�������*8�_VZ��1�*8�����ΥgC=W�C<���A�-bC�����h�#&6dٖk����.�m���_���8dGM_ʉ�r��8��R� |�αI��6#���g���$�A��y�:^ܥ�ɧDg%8
B9BA�	4�G��u}��zf������|�R��|�����2bV~Z��og8d��@g��/��(�I��yA������Pb�����%ڵ�ȭ�e��j
W�֑�P�Oco��e�o�%r��w������ά��a����T^�@a]�{O� ����;H2�=�����֚�8��r	k bן�eJ�����ۋ���j�Ӑ�uz�Yr7�$0����5�;:P+Y��h10x�>Y�R��C�|��z���҃,��x.} �C`�)�3�5�=�����ӈ���o��2]�2��Öl�5\�?1�+z�qC�C
��V)�]=��b�����l��*CU�c�SI�~��jO�mOz
��d�2�i�(�/l:��1�y'1�+Ցk�/s�g4�s�;��.TubÆ���Z�QÈ��i`�6s��狍�:���ԝsF���Ϻ��������e>!8B��΄��/�1�T�b|MB�6��p˙)Å���2ͅj�\q'p�&{�t����e��,���$DZ��	꒟���C����m}���s[3�h�Ț�ˡ�ARNr���V�q��q}���N�.�%�y�e�?]��o��c>&��Y����@���i�v��(۝3�^�(.��n�+��X|�>�4Ө��uH��,�������Uhg�h�$7����2 �}��ڴ��sr2ʹRF��lI�8Ꞵ�[��y>�v���$ÇZ!��{������!0���5�%��k#��O=�G_�K�����{2+T�m[m�n�Ù�]��y[]>��~� ��a��
Ov��yC��X�C	k��R����'W{��ޣ������W�>��X|K^�B�t�Z7	EFī[A ��+�2��2����]Nu��ɠ�mj5]a����:V�8@��1����osy��2�O1=u����m܆�g�����w ��� ƨ�5�&ej��p��?-J?o�jG	�u�GK:_mc��Cb�;L6T��唕���D�m�n�	5�o���m�PV�c�͊D%=��3&+��r��v���Q�>7���A�_B��9�U-�Š�\+5A�uy��o�Aܟ��h&{)pCX'�|͒<!�`RL{��zK7q-���-E�V&�K�[������6f����NH��F=zI������^���lx8�&��]*Ѯj+�v)�Nt�)��mQb��U�O^�r�,�|lX��0O)�+��]�)-��Q��e5�����7e��5�w\H�S|�Ы_n�
����_q4��n���1�������Ph'i�[v2���L��M�&��T��빭�"�HI�����f����>������� ������]���u/&ഉ2�^Lq$�?N�!~��E�p���w?ٚO���͗Э��)��ę�������m1M�<�9O��^�s�u[M�c�s�|~и�����^Z��f[TY�!ʠ%&�jC�0A:�k���񂻡\�V���p%^1��
�*�5���+�u�hI���1�R ����G'�V#f�n͎\ų}��wK6�T��ھ��zi�#� �_Q��J�O@���=2���G"����J�t�^��W`���5|�4�H6|�Ț�J5%R�6i?��%m�״�����lW��ڎʴGe�sT^���w������ �#L�v�s.o
��غ��3���Γ}E5}�c=��|����]x樰o�}����JtR���Z�F�վ��
��7� &\I��.�u1�uZ�S,��Ś�����f��{�O���VP�����d���v�o�P�eH4a�X<,jb�]�MZ�<��J%<���4�nR��	���?R�9Sp�eċMM�+=�;c�lsC}ݜf�`|j%�4í>Xn�e'e�
D����d<�	�@��5�Va�f1un��5��u�A�>)f�������b�+�����Dω4?\ǝ�[p�0Ow�l�	�$5��b�������͖\���r���r�r�9>�_��;�7�l������X����\��v�'P��������@I�~��+H\(��MW	oG�����{�rNt�2c�9�`ԧ���aOs�_[ij_u�c��#'j�84D"P.��'�v�V,A�h��
`�҈R&l�"o{��C�+lL����m)��[X}z}�b��C�N�8PJ�bU�_,K��m�!

�	�:�f�&eﲙ��J��.o��.��AK���;�^�[�"�LC��`�{)�N��&����sgw�\�a���ۭ.���ְ����h��YI�C��[�G^'Rk�/9�bۓ���s��.k_Hu��m;�z]?�zl(���1YgM0V�� �WSP_�sj�~��#%���E?E���vV�ǅ���y�#jg�`�o��C�hI0yL�8�����?�A>z���z8\kG��_��p($�������� i6�p�����ii�+���.=�����-|�i0�e/�i%Tg���K�'�wܖ1+��j_�I`�G�鸸�(�~������0�,+[������6�z埂�ϓlЗ�qQc��؂��S	�srK��1%�/�~gw���Q3�rrhA@\��}p�f����nwG�Ui�uM�f�E���kF�&�2���Q����b$KՌ<�QdJ�BY�U�c��ٶ�*vPۚz�� N���[�Z7�I4�AT�y]v�sz�&ݯ��-#ʁ�!��'C��%����G��	8r����T|��Ʀ4��v�D���Ϩ��m�~2~r\/��6H�l )�A*�ϥ�М1߄��/C�]�{_��H���#WS�l`��3�d��^���B�$_a�ߋ+Ȟ���npZ E�F�=�*VZϴ��nx����x�U�xI �ỵʬ�@ŝ?�b�umD��\�������ge�I"b�8���Xf�p�aM�O�ip�����?�_���	�F0�	_���|�f1d��iqn�����J�T+e���GE�� .��^3���E#� ����M,��In"
Ke��˧���rz��ݛ�m���Q,�9�bbTԜ�����&&z�F�]�+�b�g�AE1և��9���9�*/j+��]�s�B�?N���[
�_g�;�����o�GY�.�ҵZ���u�N'���F	�b��~9���lIz�L$8��3�'�v�N	���'��0K2�j ����66�ݕ��v��I='��ܯ�����J�K��8N%_&��>+ѳjM~���5>�y\@��@.ԪLKF�+�,y�Lɲ`�/p���E�p�eaНMY��M	��'Y��|��^)��r������\$�T��G^z�c���������*��S9��)K�I�6�bH�EW�,�����N��s�}���	��\&��R�P0���x��A��?��>c���dq_E݇��Y
��p3m=�L��<Ȣ���jl�?��t,`�O=r4����Hg���%7r�;s{@��s�UE���E��^�"���}@ߤ"
/b�r�Z�sg�=���1<�����b�=-���/�3$+��@��ۅȼ�[�쮊o";�/C��p�ĢA�P�7������� ��]����bB@�:��x�b�}�E����Q:9�]�mnOrZ���@�����:��	'^h�USsyN��oIFun�6��Wtz�򂺙^4wG�7�Z�N�x}�2�GW2�zw�.�����T[�8������|u]b��Qe��<ě�� `���Ռ�""��x�� P��;�MV�wؼ����#r�z�^=!�I���[A��t�o�Zg�D.��� �X��B�]�J%=�����t��
'􆽯��-Շ%��>UA�+��-���9ȳ�A\%#+9��-z+#��xė�ak�N�P�1�F_������E}� �*\���U����V����CO-js����U��>��Y�i���$�@]�a�WY؎}&~�2�~K\C���A>�o��$�WQl��E����x�}
�	ԁd��w;��Y���Өd�n��.�\�b�k"J�n��^d>ʨg�A(D���r����f�gf�'$5�)�5t"�S�M �ֺ�(���I���2Bj��ۈ�2= ?����L�5�f*��|��~�3�5a����s�S.
YK��Rq^��sQ�pY���>��IR�u!}���e樶%*��܁�d�Rv�����g��S�o���xL��08��ǚ���B�W��k��Ϲ��70�}e���cp���lFo��R�V��=o��{%�v@����j\����1�@���S˒l�6꼿	���ն>P��35sa)_G��@1��{����W�6=Q����F�^zy��&�؂���_p�=�v�?��.�#�� �wC�xt�a	� �L�/D����/�����M��;�և.3y�P���^�R�N(��_>�1���m�ў\�3����Sz�;���W�÷x4�8xZ1�S�oS�PѲ���p|�y�9
+���z���7.��a[�bOϾS_�x�[	��8��-�'�u�?�^� ��bJ�Ȁ�}P���rY�Q[оRNl�9��EH�;s�^��1�	���H�KLL8���Y�����Y>�!j��\Q͑��*��[��KP������ �^65����sl,?c�tS�+_�	$2  ,ۅwil��у�h��� ��9_�fBF�C`�!%��~d!�Ⱦ$�/��(�������1M-+y�/1Q-�4� ��ջ;�G��U�)���L%�������g����@+�V��ǝ��2xQ!L9/�����k̖������ �������k�$V�p ��ix��f<����[���֓2��۟vE����u5���_��.{7ó����	A�(y�%l�
ײ-��W����C++��N9��=S
�� ����������Qms��M�����#V�?bY"��n�ȇ���1�w��o�{�&��~Ű5����H���q U#_8t�R�2��~��Ѷ�r��6K��{ɩ�#Oh����p�c̨�qc�eKe��� 3�;H��̡lY��o⇠����ſ���$�@u��Zu��GU�ˇ���dGE�6?B��K��[�T��G_��I���sʠ@e|g���u\4 �q4�5��������
<�������lp�Kې�B2>�]�c��:� dS�l��X�M�ֹ���Ox�N��[�;���P���8%?���T�l�jw��`��ξ��Ԝ��X���?t������9�<!��V����������?g=�y�F��d��}�~o��O�"�C�u����*���̃�+9�/rN$C�bA��X�U�>�ٶ�Y�K�K&������P�r��S�4^���Ko�z!Lv��%G�җ��Շ_oLq�FpY�P,qN�w	=�爃���J��\x���Ӂ4gz�dT�!�t��#v�V� 9%-Y�m�C�X�l���Qc.�~j���/FYE��`�
��k��
V�*����B��r��Q��A����)�i���A�o��/%*@M�0e���w����Ġ�\�oN��2J�{Zƀ�ؚ*�x�Z+��Ƕ���yl-����K,�C�o�nZ;�-����TK��nW3��3C��:�R��A&��������Xra;6hS�(�Y�!	�;l�M\ƙ)������@m���%�tM&L�׾:/�5dp���c����x���6+�����C���L�"]D��3�p���
�xHʰ�a���k��C��F*zWcvB�"�5WKC�?v�w.�����a⠧�rj���st8�Y�q!�;:F�9��j��!$��g/8n@=��r(k���c�_:ÐodnW� ؚ�+��De1~�0n�?Lˈ������G�m��l���A���ufC�(@h٫��ٓǇ�{�_�$�-��&#b��<<zW�7=�l��`��&�W��Y~l]\%�\JfOuQc�����H���Y�:��~�f���7Z�%7�|�N���x�#hr�0�t�;�:݊�þ�r���u��3� �āb��J;d؇c��Xj�)�;��E�:��Y!�#�Z�-f��{Yv%M��]�=�.�����I>�(�+���+'�҆�n%ˊ�t��P	y��&��¶�!UT05�Ԃ�l�YC[������*8�� �#Hm򌋟6^ �K������]�+�z����;�E�.C�Wa���m�E�S �)>h�.$K�Mf`Ft%��E	1��wc}]���ΆTVh���E"N�(���X��Αmy��*8���]@���[7C���ń��Ce��S
a`[@�)�� ��Eu�I,2�\k��Y%�y��{bA�$�8���H�g�%��!�Q�˦�%WM��fpl�\�`��E{��j�W�h溊+������f)l�V�L��j11W�q��e�W~Ҥ�^�	�s�̉�X��MF=�n�B�f-���DO�S�iX�P�p��=X}�r��p"���(FU�[�;����ٍ,��7¾/!��=�kK�x`>r��S�  �|�瀕#kǓ̲�oQ�>��/Dh�D�v����U��d(��/��ҭ�P�~g�17�cQ�����P���#h�J#B4�r��Xa�B��s'�tIeUk%����Ӷe�PZ8g0ZU�D�ۇ���r��i~�8tvk,��Y�QF�Bff�7�J4TB��N0�2�S|Sr�� 
�4.Y�"���%�^��$v��X�y8�X9��e�ْ;!�vZj�)p������9Xa�d�\f�����:���n0).L�,��f�KC��1�@�k��Z%�_y�����̐0{/�O@	T̕�ߑi�7�ܔ+�>���%Œ��x�Y6�Wd�o���wΤt�+�&5��?�^�p�6E��8�ۀ��rh���E��D�T]��Z���_���J��(�U�`����漶H�B1T_\�wĲ��V�x�����5��El��j$�#0J�);-�I�i"��� �z	�;&���aY�:_��כ�]�ӥ��ɯ�tJ.o1�q��Tu�;��F`ޏabߖor���L��P�;��#E��%+

a�ܑ��O��!g���Rkb��dzY����v����)��@��]�":+�I1��H2�*�>�5��A~PPqM��n���ΰ��s/�M��MF��8*?�aݠ�� �"=������j�6���	���k�VoF�~z�y���w�c|$�����Aҷ'`08�>+�1i��~e�@��q_�|�E�j�9LP����=q$�� >�PD�\�W����f��0���MA\�`^�� Mb��[O� �0��b �ak꒷0K�y��o^5(U�����s�=yIP�z�S�^���{^��n�����"^�7<ݔGB2k"�@xN����Nq�g�%�mu���d���9G$^8����8�)�3d<U�Ό%
��	'!�A+C��
=�dR�ω4:�S���Ӻ��zA�y��/�,�}�j�GuM"��eHT;u�+A;0[9�D�ۣ��?Q$��1�
�>d�L@_1����.+W�"��ra��^gV�x���?�����|CW����s�J�N���R!_� j���~9v;�ۏ�� �Ʉh��ރ�"M$MW����8wn��2�K���d�}b�}$ײDf�����¢�������I٤��-�\k���
�`�Z�I��A�>Z`�0�u��@W�c���$�d��h�.ҏ܎>�5�l�Z�ӱ�/����*����Չ�AU��ӷ!qQji��n~�.8���g�-}7f�u����Ɣnj~a���6���}�mL�=��^�����q��8��ٛ�
Ϻ�|�^�l��B�xwnM�D���own�<5=o�!��`�KE�6j�����i&jp"�{tpFQ"���ק�%���5�wN�]��u�Z�����ϖ.��cx��~E�q��@�@�,��7��'}��7v�q�xъ�	�Ѓ!��?_q��;�%p�5�=%3��c:Ɵiv��7���LM�^Ą<-��_���f��(��fʥl�[�^���F��tћh<�Te�<��b:+���t���!+I&��<r�'m�� `�ҭa]�hKG���hx;!��*��ӊ"���0�L��i����Y�HDm�K��
;�#����+� F�,6�DE^-2(����?J֢Ī�:�D�N�I��%T��b�Q�L��:�2��`�a�|*��DZ[?��<V��W�[�y�N"y�4Uy��҄+?'�5\�A�7%�7�P�#��Qn!�L���X5��ń�nS��O�v9��@���e� �%i��O����MuIc����]?��[�@`%#Ȍ�'����2����L>Y5|Ž���ͱ\��d���c3&���#q�˺UZ�cb�*=Jzh��\(�N��,	8��`Xt����ǔT ܇�*~�O/|�2H�HV��_�ښ�7Η&��u�{��0=L60*�T�p����_�K�LH�� �0��7>L�����*��@lV���Qԟ��l��i������HJ���G�`nf���E��?h�5Yu�����{.�Y��I��#�5lM}���zg��n�y�,�H��Ce�<�}ZZT(Q�Mb���_Kс~>�����^��smܬ�����o�~Vs�`nY��! 	N�`�'\O�p:�4Ǔ�������Z���+���P����y�i�
WܑthTS}3����w!����⊧��G��L���=�Sς	&g��C��C������ԟ��P���!N��4d���:�/�t����'��*Ntvu�c#�(;z>f�|���kb�⦕�Tހ���>��.5��	���L�qٗC7ဪ�P
�q��<�
�/U?f�&�|/w�p;I��9���g(���P@S;�6��D��_ܟ�ԏs:a��a�6*��ު�w�̶�����;P	��#9ʸ����H�v[/���<�F>4ʨ(�\4���.���w�Z:�#��6̘��"���M����B.��P����Ein�3A}�'��7�:1������:����:���-C7TW�E��}N��8�X�Uȁ�!���k:8���?��Ե��& {�(���|`�<k�Br9�i�h_���/�!��l�����o�ps�&!y8+��F=/6��"�](�3�����z^놡�nA�b��߇#��+�{��l�@'�dǄЛ:́L��]�ΞY~����/�͐+���Ĥ�x�DV[KT"0d6�����@6{�M3�2l6����cqS,,[��U�o`��4�������xq�ӂ*��Xs��=��vQ��OmY~u+s�*���;��)ɣ�����?���S�b �X���p��С��g�l΁�x䨁�*�Z�K��M�,�i�+��f��C.鎰�65��,������I�mXd����?1��~>�w5�A�m�!T�k]��ޭ$��2����uI�F�se2�\�����cH�R��P�,\�
T���HW��zl�6����eeO��N��и�l���~ۯ�˴��I��ꎴ��L�-��T`,잖0v�r���@Z��`)�)T�����,��Z��+���5�ŝ#f7G�S��w|��:[��e*�K���h�%8�8�;���H�Ŏ�{������p㗆�ۖZ+x˫�SȻ���v��6l����mu��q�����ܴ����$�#J0�P&Pe���/��m����Ġ�
& ���k1^��5��� K��q����h5���8�v�jC�6*�
hv�m�4�	T��j�6(����fޔ��ƙ?������$����M���Oz�'R� ��?3�ر��g(�V��o�o	���P�Pn�@m-����PO���9Μth6t��Ti���,HZF�oY��u{��6�Q+��#���D��q��Q�rO��!KU�dc�3|KG��Y���;��7�L=f�y*����)�}")��.�p�s ���V��u~V���8}��?�ڟ寺O�0��mYA�5�	���� �j�?��� s���0�`��^��q��J7a��2����P~��AfT8��g���Q���@�!����LoWQY@�Y*�[I�{+=ֻ�{&=,X���"��@`����ز'�z�r��%�"��t��;zNUlf�g�o�	B�qf�$xl���A)p��٧�o��R�@��!a�I��e?�N�v���D�C�Ʌ���#B�~�Gp5��qO%Uo\Q.�>��'u�`?6�[�l���ګXopY�/������sr�Sg1:Zx�8���XrG'����@��P�@�xF���v�������V
h�%�ͮ��(_vS`H�2-K��Hd�t�
\ڧ���x�&Č�
d�X�p��!y��Ĳ��cK�Y楄����!����Ux�
�m��� sZ���2��e�/7#�<��)�+H�S�LN	8���R���7��'�B��18Y��ɴ��_�2Ēj��'.a����1e�K�V�/���彦ܩ���wE��X"�X��{��
3N7���Gj/?�E1�b|:fs}��h�����cݠ��xu0��a'H�M̦nM!�u�-l|&���D�#��w���<�A��¢���)N��تO�g�?S��K5����1I��J����(��mo�w�?K��
>���^#�y��;̞�W1z���T�{��|���Z��]�1Y!4�[2�l@��*C����	��Q��T���Q"��{J���f7\k���k�Tk�悔��,�d��R�ʀ���4݄_�es��oYGDN���ʭ���F���?<���[�FX�7;+IxL���j.T��m�CJV�������S����U��i�y���U�]�m��,��h�yUxX�I��eW�����<Z�aZ6�lk���od�Z�凙X����$$��p-r�B]<g@�%_'m�!�Ik.�3�{uph��éa'�b!"Q����r/2�%�\|�V}".�� O�x?�s�R�DΖb޾f�I�~��мRGlz�y%A�R7�G��I�S��2����T��*B(�y�˅�ī5���KJԎ�==|Gl��n�q*��b��F?��9��g�f=a ��Z-�������&��\��f��s$�3���d��<����X����j�О粡^�X�X�+�Ԓ7�pD��c������]9���z������s��?K��\�lxi�#y��֦t=�!7��H ��s-�x{CC,�X*����(���<+Q��:�v+X� ֡z��L�
�	�WF@��+��*B/�|��G�r(��1Í���	��7W"�'�ؗ��Nyl��_Vp���d�]W��O��<COn��DG�Y8ωt}Y<�b{�ș�6��4�-�R�o�ە-x2��:s��6�4�Y�?�ȭ^�zyftA��G���d�D��S���%ڰHQ=�o�rA)H���$�k|��a

!���|%G��&��Қ>�V)�r ��
̥؋邂p���n�h�p�h� �lrT�5 ��7�;;1��YU�n+;�cq��X��C�&�5,}եc�2�G̬�� yƱ+0�p�^(����=
�f��wnG�e�B#_P
�{z�ڤ�Z�Jv�B`�y	�'^Q;�%�5ް,T*��%�h�(X\j\X�#s�n3������C�$��?�������������A�y�ĵw�@�35�	#n�������_MM������NŚ���ՠ�\��!����Q��dT�>�z�@�L�y�`�`^[t#ϒ�@��/rs8<���Eġ'w\:hi(��dw�țc��rX�'2�ݶiA�j6ao� w����v$�>dm���\)	D�� ݗ������B�z��6��N|\t�q���Q�۽k����t�#ok!m�wLqr�'�7����U9���
������kl��%�j���s�s�m�_������{��x�b����1��]�ej�q��XeK8�RΠ �����|�9����9�VH�����+(5��`|��U��W�<B�7P����PO���L,���U����1�}�n�vY߬�� ��u�p���Aa�5���SVat�0
�E�����.�J#R{�b�j,d���0�Ѳ�����kGh� j�-sc ..�Ć�����4�~�^z���J���r��v����M�!Ei�zo���g����C��좝V1 �)(5��onÑ�p�'������熠�����<��It@�'��ˈCY��Yf�1��aM�.���l��#�������(�>�r�P��ۣύ?	���e��L~ph�߳����(�[�"p<�9�-|}e��s��������^���b��t�b�s*�]\n��!���eZ�g�b}��43X���:�s�G��H�f���ߜ5K1b��2Y���-Z��t�	G��j��O����'���N�7�䵬E�#{��ֆz3��9��>���Nbh85�E��֬ ������O�	���-��u7]m�i�M[�WxL�ҍ��@�q�7U�F��_;^���oY�K�r���;���-���P1R���BP�#DЁ��Q�����&T��*BmFqJ�́��/銅�)j�^�`��������n?�Y^���
PbE��v�p\�/<�o`ʴ�+s�VTE<i�ʺ���X�-IwF�^�����E#�����}I~�.��bJ��I�/�b�}�oV5c��P-UQn��V�*��n]��Z�%�s�s�y�H��6��Kh@�N�G _J�s�&���,�A�e�l�� �[��ol%�ZK��Ke�s:ώ��PV+H������Ůy}�Yջ~1B9
����>�9d.��^�;����`Y� X�W!T�G�,f��4�6��~uoc���X��Q�u�>��>��N`:nߒ���]�&ꂷ���x���[N��V�����( x�τb�(F�V�X&��r$�G��2�\4 ��lp"���LQ8꾇���ۈ�)��*�j���r_�?j��㢉�q|����<,
\ƵX��奎Ą�����e���r�\�ȭ*��K)���b�[��ó$"W�N�9�.	���YQ�v�%��}���P�p���3��+e:��xn>hN\ˣ� ��ù���D��ȋ��RIuY2�t�F4���)J����"ښ���G������ugʤ����y�c�+��(�u���V?�U.!*f�\�Q��C���IL�R�p�	�z�[gmuj:�ۮ-nhp�ڑ�t���B��B�!A���86ZL����V!�z���EZ��"��ݑ�ů�t�>�9����b,.[2���b�_Q�U��b�"!���G�e�An�Ye!�r�q�fO����P�H��a��;���S��~�'�L���OK_AMe��������^aV�6���'%�_�i�2`ѿXrEr��<�@�x#�������:��%[�/6]���+�I�$l���7���;�I��m�d���V{�s����zFa��!� j{���{;�c�F P۽� ���X6P
yJ˻��wE��Zo�MwҰ(1۩�+��<]pxmi�	?��s��d�4�lG�ؿ�i��u����g����'���8��4��rˌg��{�0�8^������-/�I���w��4�@������[u��mCܻ�t;���i4��F)U��Y�=?�Z��H��E�������f'k��q(�s�ߑ��;��]u�aa�\a΍�Dk��~����*�[���
�sw1Dd���E������NGO��
㌞�ظ��D,鞨[Ր^@^�񢧮�ƗѰk������쳞���m��C=����@��������P2�湈�_7���E��_5��M�m�y�hC������/9��*���[q�ݪ
���]G'��xE:n���j�.r������=;���ҤV�/�
����P�Yc̕a�E��#��64� ��ǯ����+SE�Z�Ԍ
�_�W�j˸��� �F��q]^���1C���s ͞�s#}/omVT=VP�*�]L^)�b����%�Cv�s�Wׅ!`����^{y�_�n2�*�������Ӗ�S���d�{�������]�ah�����t�l�/8��@�4%ĉ$�A|hK]��}��E���9np�����%�d��uZ���}<f6j����#�������<���Bat��O��N����4�n�;"L3`� ���މ��@��s���uuۋ�� �!�Ԫt6~�;��R��+�����w�5�=UA;A��r_�z� <�������+�du��W���9h�z=��� �ᒧ�2�]�e�a'����p�V��=Z������N�/��E�t��
���l��X b�֞ sV�9T��5�,���J��լc�(,��9uE�^�b�VA�Wv���sW���6p�b|:�#Uv��
HX`
Zi���h�{��'J,�.���^��e͚������_��������z�����5�RyRŞ��!��v@��@x��4���ܒS^Y���12�Г=�F�䕯X�c���*B��Aa��9%3���˜�R1�z���Ha/��?5�j��hR�ڠ�~�~�^���$���|.��T��^�������w34TU��v~
?3�#�B;9�F@�U�KH���*�3��͛�u���AU���5r-�4Va�v���9ؤ��,��o|�a�mC.�ζ��pׁ�"�uM�[�t�%��wt�?��4��w[�Y��L�=v�$�T/P���c���ޔN��x�J�Y�BY�ux��g�o9�Prҟ�7���c��r3Ő�@�b�8O9�P)�םb�< zj��4�޹ReܼR}�A�p�5��������閬�嘩��9��g 7.jmu�6b�r���B���N]j����&�z��Tv�9��۹<����B��VJ/���R[W؎�����0�V����)�|�=v@Z7M6�֬�V��9.���392}B:��Oc	,�U���K�@��^����~����Ԑu@��
�9��ei`�x�D��fNV ��sd)����D�B��?��d�şQҦ��6�5�۝�Y+� ��/�xw�!���h˚mѱT�b�K�������!�����k�n̘K,��������zƕ,��a�4��xc�l���Rǆ[=\G�_��|�x�8!-�л$��AuL�w?yzd @�����2دT���rU��a��]�^W���b��� b�!��4V��<���D��צ����E�����v��Kd��Ѹ��!꓾F�vy��yn@j�G�!	WJa����"�h�[��'l
a	C�r�yX�w���Q�^��B�"��`��R�$��[;�C@�;�Kc����Jǀ��v� �S'6p-,����Q��A'{V^	��X���1�>D&��g��#�M~*k�پ���#[��R�B�eb�+c�����I�Un{I�ʍ+˓텙����L�N�� �-��`b���&�7!���\������:/`}�f�h��/��ߊ�%�v�rA�~в��Gz���#._`Qu�J.������`���$vg6��GY >٦c5f}��z�,A���6�z[��Kc, �3��X"�KP|����F�R']�I{5W�r�u1>�4�E�?�{ ��=����-6{'W�Va�o02Q�.ǚ�W�T�3�r7��o�j�.%ch�U��^M�����u����5��P�C�O����6b�lC��-�B�G�X��d�ɀ��R��Na-T�)�+�f����Cޖ�z4�$��y�b�S]_���<3�S�v�2��f4~���0���b�E��cr���~lV��д�&MI�tK,w�	�o^D�5�d�Wڋ��;z}�V�r��șA!�bz��:��Ud)C�۞�ɱ���B��ݲT6r���(�f�[�PDڵAg�/�0A����u����_<���Q��d�����U�?��Cܮ�Ɣ���V�|�1]*�g5�X�|�dcP�;㘾>����/���|C>��gI,
��� ��M�����Co�D�N=0n\�'Q��G��'6�C�a�|��A�e��M��?e��N�����O�<%R����ψ��Z�\>ؼ��a��#Y�7�݉���H��J�,8�2���*��u���X� �%�^�j�����$_�e�X:��g��EF�B3+M.-�4J�:B* ���\��c٤Hm���GN\��xzs��G�F�	w��_捎�u��аg�|�儲��d��;��"or^�`F�l��:�UUϥ����J2��hN��_3�-�3(�D��oE���ߪ�I�8�n�7�CJ4:�h�P/�5��]���S�t��`͍r2��3fޝ�"��-:�8��ZY�@7����w�U �o���Ϙ�kiwU8��$>�,]D�o�{2	|�:�n�|e���p,��k�@?U�4��32�<W��m2��xQ�|q���eӭ���E'V����dN�8e&�j�)��e����sG�+s��nL=Ek�p '7�����\��9�UV����Pn�Α��\�+���9�ȡ)YF9�u�ݘ4C�XZ*�����n����z��-�n����z�3�I�"n���P5t����}��(����--%��g�7�Z^*��HK��NX�G !RP��%�5���9��2�܃�JC�M��i�G�R�di��{i���FWhHN��<�5������a�3лQ2&���]i�أ��9�iSFȓ�ɇ����i���!�����g"e\������ �G�ś�e~�u#�RX�m�Ȓ:|����Z߹�9;\?YYzu_�����W�})�,�\`|9��I�K˝�.�߹_�}�ֵp��N �^�L�Sr�	8 :18���Dl/�0���u��d�_�g�3k��'h��t:�l�0����IǠY��FI�����pШGA�i� lDLܫ
Jݼ�$��W�����0�}mj�X�M��ٰD�v�*_�;yo��w&M�<��:6�����$(ׅ��_q����Y��oU�X&瓽.��@\�3��7���sQ7��a�ł�a����r��\�׊�$��������'�Y���a���e]
�q��9���8P����2�Y2�6����L���۔.-�
�gw�rm"Ų@O�� Ȧ�l�4�<H�@7Z� �����T �'����׉�
�(s�?f�@L�T�|d��G§��ps�:�GNBT�#n�'�5N�_����!hRƼ�cX�ry�5q�VƊ���~�"GS)������ ҽ�?vݠ�4�μRt�fAXu�1��!m����fQ��l#��K�	Z'k����X�ʈ��Cr4����:4.�_����
m��SƋL��9U�m�Vf�WغG��F�&ʧ^/�h� ��ZQ��pN�$�E&�7R1�+qd&���2�\����\|O��RL0l��ಎɳ��x�Q���%���c�n��Ҹ[]x��GD�"R�CPmU-%�^���*�
��4�H�.��Q"�6D��
�>��v�ޖ����Pe�<4�C�Y@��7�7�<l��uޯq�V	ć�7G�t����ٵ/T��W�S�X�	Ҿ\���_�V����nM�$�m�<=���'#3�D��D�l��Lj�$���Ԑ����:]X��&J� a �.��m]6�N��g�,C������]i�C~����Պr��Z�R�y��ĸj
�c��g?���Nx؜D	�~�e[���wm/�&��R�؉@$V��@��!�T�$�&褐���	�"��%::��M���p���L�����קd�4Pj�H��eXx�U���HZ��/<Sx��@r����	��<�iW�<z�ѳ����Kg��y`;|��,�"��+��%��c�����X�5v�|HK
}l���S��nK�l$����"T���-KE�x���>�+wǩ.��3\]5l�X���� "�����ߜ��aaImE"�6φߧȝ� Q�Wm��y�e3C�Ã��'�b�@�E�����lj|;����y*Pz�76�	nD��'�XP��/;�V���gO.`k4���K��;4�hŤ����`P�&�o�8�g���4���/O�`U2î�nKK�����C�R�ň	��1���N�<ܗY�H��4W�NT��|�'���9��������������Lդl��1�)#|�=[/����HO�����h/��z��g��O�|�'ҹ��w=�8���V�@�X�Uu�q�m�x�	!�8ӻoӈ��/r�{��8@+��%nvH;����rz��5y+�ܰ���5Ѧ
�k}��OW1�5L"�rW�U�=�l (��s�ޑ��R�J+q7x��֕���Ȅ�m��|ݴ�*Bm��6��M������yXa��pC޺3�i�wL ���7h�X��I�򖬎��1��?(j�
%��Ds�C�Fe/���8�E]��&1�Z&��֪�h.�it�]ߊ�`��C��Id����%����{�I�~�aNCЌ���s�'#g=�}OC����ӪD��͢�������8:z��E��/o�Z�P7I~�� _]�~4��~��'r���Z��g�!��;�:��_._��Wh�[���3�
I�"i�zjʞX=f�)/��Tmb��Q);ο��v+����㨀��A��Cu��G���)�<!�׆�i,��+y��f�����<&M�g�x1�����m���MV_�덕i��r6��ӽv�|\6�#�8х��}߹/� �ǟ���*&�]6��k`&��D��*FoD��@��R	��{�����W�A� �����/�)i_� d��3]�yßѩPԛƆ��(�?9�-�f�*�!��\��<xMφP�̶yeF���E��2~��7����w�F�I-�|r钶O,g!|:U�}���\���wd�U��x���U���4t�_���ҵ�N�0Ź))�lc	Yjʦ�[#ϩ�1ի��[���pt�;���@����?����h}�Rv���C�VQ�cۙ��Nb���K���MX�����U�uR���W�>̘%&�%��3>đ�!�+h�qn��3�0D?�0����[h<�|5�i�		��F�d��y���O���2c�����0)]o@g�:�s:��۔=�=��Iw���[N;U����[�b��P��kk�h;e��3V�ok��;�mU�M�U ��Fҫ�]�d�4��b�)�9�S�4�e�~,���=l�ܒl�<��I����8A�)E�o��w���"р�HJ�9pV}.�������h>"�z7�w7.�4���m�o#�Y@���%#�����]�%��3�����)B8��l�>� ڛ�yH�$K�@�r�_��^~2�t7���?{��?�97 �* }��0n$�F�GJm$��~��DM�*}�P~S��8�j9(�]Kݤ���&8��'�UB\�����x��~�����B�n��J��x2�j�R�ǼxJ@K~�|3Ȃ@AH<v)KX��Up�D�gy�����+_X.c��ۧo&��S��+iл��}���u��K9�T�Tq>��?�=CVQ
�Nn�{]���za��%�Xp�i��'�~/|���*cm@hrb ���z́�K�YD���W������;��\�ڏ��8=]����{�\���u�m�]Y��s��t]�^�f�Iv������ �'�3��c L8,����i��|��C)�8�?�	9��@���|���@�ׅ��?,o�Á��J#��@M��Ŭ\L��d�أ�Şo��jy��{ ]�?$��ʻ�B�&�CDH����8�
�05�R�3���%�p���2�S섘�G5SZ���r&q�u��>v(;�J��x���9����^|?�؅�1�!���[��߬���V��n�`��v����!�Yî��������O�C&��kE��q6χk� <c�2��%����229Q>����c�}Y�*O�h�dn����\�Y!�fU����dM%;=w&Q�)K��v]��b�����.�	�n%]o�,t�'ÞAS������p��,�����"5�$����PA*sdO����S�3-=��?��Mc��E	�G?�ZR� �t� ����e��0�bS�TE��_�#�{Zqdg�o;�7��	+J!�jc�X~qԒ�9wuHs�Y;W�x���#��"R�u�k���$^=h��䷥��U~�nal#�6�uG�0ɡ}���CD�E��ZN���q,�L�T�h���gV�}��2na��0)%7dnk�$$��o$;��a�΀�u���F�0��NA���l��9s�>HE=��|؂HVK[Pu�/$���v�s����%2TT?���&�.d�� #i�@�h�#*����8��' �U��c�^�<W����h�Q���@��dU��
���4쨄iǜ��)�n�!�nj���	�`<���s3fO����]E@Cid��M��G��ɸ�"���l?T%ʯ~L�'.v��Cm_�+� +�@��3~�_2r#
��Ϥ�w��&C�P��	�_�'��63	.r�����w�W�gy��˘*�G�����9vi�����ZzϾ\%�6����P�G��.x�