��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj;�:��H��`��e���f=?F�]��Ƥ,�F9"��FS
�[��G�aT6E7{$n*��sS^�3�B�؉ҕ�1���<�b"���2b낣Ҕ
x?�&%dJ�8L����$+y3�D0wJ�| |ͽ�yj��U��r�R���Q��muH���]߿�XJن�3-M�
�,��W��ެ�X�C�;!�u���Nm����S׻|��]:w�.�K�Q�?2^�/����X�bj	(}�wSF��xIFP���)�y���V�RL�V����N�5���L����  �H�=��J�"�(���\�'t��I�tm�^���%�iO@7��<i����yJI��+�߭�z���������'�"7��U.M~�}r+2h�=��YF.P1rI�O��8�z�CBN���֎���1<嵵�aN,nVF��+��}v�
Z����8ϒ��B;���Mr����s�[���O_�����H�="$���J+�).�zt/��7~ �m���[��P�R[Gw��}j��s��E'\L��pR���e��s�`|�,
�:��_/x�:��T=����'�Q�z��[���0}���xM�Z���s���β���1��"ں��S�\-�'�g�h��+�7M��-���H0�k���5� r��0&EL�<܌S k�n^�L��u��� nNv�BR�����<��ׅ����1f�%X���+gʏ�n��i��iU{��A�ڐ,��ThO����9�,��n���b�_;
+0vz��C�R�cߌa8��@=����K�{
<��w�"h���6@�{�[�����[�f�v�v��(R�#3E��B��9��YV�2��т���!��8Q�a�-�M�b������IC����j�p�0%�b��s��-2�	,�����d�"���|/��UR�15]��nL��U.�F?�X���D0c? �l\h֚���f뷢Z(��X	0W8��){H)���K��	�*��J�c|Pw[Ŷ9X���"wX���6h�X�Mø6���x�|��<1��Do!/�J-*�,_���Q:j�qSLA/B��Zqgc<��> ��Z�fy��Zs)�j2V�����9��	�7V=�`��Ͼ���:}'�&�r(��zx���vӃM��&�m��l�&̷g}���Y�͸3דH��4@~{17��E���dұ�3}�xZ���/�]�?�˒i=��!����I���R²&&�� )34����F���HMX
Ӯ�ˬ/6���i�}�b��x�n�q�X���ݝ��S�K=�p6�Z�m���#0���sя�q��_��4�{3#��H|f���q�1����)s�^�N�B�ߞ�"�(�aӽsD���8I�*W��ph�-~A4zr;�Ք���[�$�T��\��	�RȡAH�Hm�S,=��n]o�����T+A�j�ZUWdqXJQ���8sܶ]H��7��mX���F)ô�����q0�u�&r܄@1=�	i�~M��!��J�U,�Kg�~�W۔�jq#=b�Xs 4�"5	�u���7��Jt�� �ԉ�O��ޥ[G��
I.�{eJu]5�g׽|	��Q���,��4+H~�!��Ad��ᬲ��n� /����l�n�8mj�D��V4���1�3.�38��v�X#�`�K��p-�b%J��MmN����Bԉ�%3}_�-��tА	$�9�U� 8Ƃg���0��N�6�����4Й�Fw[��:�qK�dx"¶XW��K�d1Z��(�ښ���gs[!XF�{4��_*�kh
�L#ĄK��&�?�����@j��DBr�.L��&�]����0���[n��Q?ϭDy�t�lg{���_[�oCjbK�u�t�����=��^��G����#�8�2,�Wm��4��eӬ��G�.�I���tbԵ(-"��log��v�ƻy�}}���#�}p���F�/�7�F����R�?%\��Z�O	�>��>����p�T��2A�/��_�AH "x���N`���بTr�;�����C���lg\��eR4V*⬻g�#�M�[�׹A��%���]��V��>�=��u� ���e�ފ�^n~���3�QT�IW2�y���wn�3$R�P�1���؃�m;�~�ɕ�}�n_���\����f8|�qh����H�h@��}����~�"=�y��e��n����"� f�ɸ���M�xE7]�(�4��巚"l��N�&�$��)[�*���C�uk�k6��<�|){G��������r�lu�-�j�ycZ� �i��1�̿�\�[/<����Kp���D�@�6�m����0��Q�MV�B(=u���#�y/�'��D��p�Xn��2��k�f�~�Y��g�A+��7�oٔ��L�PP5�9���g��{#�Z��)��%�d�:=��jH4�G��S?��@��@��g�H6Ho��Xh�5-�cYn:�7�|/'\˄�8�+$-5���(u���^ʮ1��7_"��!�A:�mҜ�0r���h�<��}b���`VI�>�&߶q�M+��Qlڥ޿��;��hjB�q���gP#���N[l֕�D2��أݶ��;���ٞ,
��{'��r/D^E/A>��i�Y�^O���?*��N��-���F���g��,Ժ#��������u���pR��=��`�6x<!b�:��"U�$;RC��y4�ssuC���x�6X.Z9�b�Ʃ�:uV��.�2�H�M^�Z�n+�]�� 7�c[wύ��>��[	�^�|�mуI/����~H#=!Ϥ#��ׯ�A��1����y�7ϰ������b�3��Fj�o�\��/�g��67�P>6^�.!-��/�؝ϑZ2��}ㅺZU�7�b��-㏎�޹6�׳�u]5ɲH;��;����X��W1 ��Y\��'����F�Y�!'v�F��DS/�{T�t)��'R��WEA�Lu�׫��k8�������A�����v��b��M��5m���T��i���A�E\��G��;t���c�x��4����f�4 ��+1�5X5-�K�SJ���|k�|d�Ͳ�������Gt[�>
�'���Ð1���
�1THN*X��.� M�Y��E���k��m��İ�Qs�Tt��ج 6D�ݼ�D��F�<���h�J���"�#F�ܖu�������3-�$+�"xq�q8�dq�2����)~�bz�5e��$����ԋi��SD��6���8���4>�݅d��g�B� òx�~j� ���2�+n����4��}0�([2L�M��e|D��zR�Ï�.Jtxt4�Je����� 6+5��Pkl]���.VT���;_ř����b���_�t�s���{6���1���`�&�,��+g�X����h;�W=n��}��Iq�?�e����|X0Eq�����I�����i�^�Se�ϸR�{�>4r��rǴ�#v�j&A�@K�~7E/ֹ��A� ����s:�<�K�G�~���w�olZUˍ��$g�DKl�ȔN�:��� ��0H� ~>q9rbvj.[�	����x;z��a����
�D��L*E�Q���� 7C��_]���X0�K�s������)��C�w7nOk�F�F��?q�a*lv{H����3.�\��5:Ө�L�-�^�+���7�ږ
�_���h>.n̉Mx���U�AwWi�/e�\�z���`
��.�y���&��X6�� �-,�ϞN����U�޶���1d���8�������T�w9��#6�����"���P�:j�E]O��&���ѫ�v�0���8ĭJ��XNǴQOVi��B�� W�c�`C�s�ԕFˡx���5^�]x�H�q��/A���e�7�Y��C��(�|KSD�u����g"Y����"f�(��;F���Vt��Ƃ�l�|J+���M҃}���>X�[��X,�jl��'�z�sy�ll��)�6p�����p�:G\�����]���rb��I���k-�UmOhӒ\#5o�g-��VÕ��y��b�}�&?���ӯ���f�ݤ�I�z�������i�蹷�0M:ZPiF���vVR�D�;W���2��.>+̪�ۄN�x��r��1�$A���-&��VQL܊�d?79' �9�} wI���E��&�`�-�_q���`5���8��/?쌦(�kH�Tj����6�G�?�[+Ay�j�i9˘�ƹLs���dqhXVf����� ��8�n�V�~��HC�?J�o3�����Kc=*���Y����b����kq4��{�x�7hG��M�F^rtO���`l InL�LE�oC���-FpiR�}s�QluZ���mO���{�ۗN���~���YC���\}A�믖a/���i#�v��Q�ʻu�DH#��H��4�r�	�ʔ�� �²`�Ld��xV��8��� }���)̒�i�PW��s��Llx��^�f�k�wr��;U�I}-i�&�*Kz�����R#��JO���5z����'b��_��QJy��p��\�V�L��D���6cTcn��|7��MB��ZA\=�����,�h9��K�><���>L���tN.��iY�~���A�=��� 6�!; `ȧơ�EV��4#���#,���	��v���3AdHUX���|Z�x�];&�P��sΛH�+td]�^{=�4 �&rVX�H<�}G���J��0-�8Q��:��S����&Z9�n/|�` �f�؈Řr�+k�����;7�bv�h�Q�%ȱ5m�;l��O�b���t��*!��+" �^���ئ0"��>u�3`v��������y�L�F��FO� ��w�*N�`�?D�6�)8���	k�ޘScO�x2ؑ}��dU!"����̯�)(c�<^a�27��(0y���yOo8E�6�e�gh�o�$6��?^�[6��b��
DsT�/���u�)t���Ӣ�ҍ���2���J�ɒ�Yq f1��_z��g)J���7h1k>�>++�,dĞ���>�S���V���')���8�wC��̮�J_� C�\0�P@wUZ ���a3Ot5$��[����Ziz�	�#Ǥ��|ϩO�j��~βE|��h��)#�Q��L**�4I�Wmj�fm���=P¢�lu�F�Ba���"�Ef�K�M!�����CYH���y�R��Q�p̂Ҡ��5��B�YY����s�[!��EU���+eL��9���Q�k� Ҿ��aZ�S����o���'��c�õs��� �I4{\�S�.鿼mp��7��2�D#����7��z��[�u��!��zM�O����Ɏ���9��-�\���I"s��'6"ʆ�,���FaZ������������6�Sj�L�������5
G���K��d)����FW�!C�����z���(5�*�
F��mנ�_�X�����%8�Y�쀔�u�{*x���2��C�r0�����O����)_ޥ��2�O��_�x{;��J�ω)0񕟞�9@�Lk���?�n��2�r氱�_��0u���x�
����6d��ٯ�Gd��ab%��Qt�H����L�����ζc$�'eS�I$s&)y��h�w쐉�~�P�X���T9I�=������M�'!��)%9�{.#>U���Zm8?pD��MX��z�溗?.3	����b����ȥ8�4�^�q�|-
 W�y7��gҋ�������!��e΂��3��ie����+0�����<�� ����o����j���$qc�d��7�R��٤��>h�R�6��$b��}{:���l�P��χ��=e⇒_0m���h�@��:r�Ԅ�)�)6��U\8m��v
R���a��?�C�6eh.��i�\hE*i����d�9g��-X1Gvz&��%)���.�V��&�K�s0�:w��DA:��7>�A� �됅,�P��||o��s����������@�%��cL���ؙ&�Z�}��H�E B���Lg���}NgUN�3�tp�=w
�2W�IˌN���k4W�JZ �h�Go)e�'�Vr}kT��ֹ8�lC p=Q6׊���mx����5��$P���,��/�+���F[Aɩ�AS��o��V�J�_��7�/��:��J v˯6���{��\�'ܤ����m�J���L�D�.��y�H+�+ļ�ů��oMn��'�gM�5r`g���	c�I�]M��d�/���a��a���)��K��DaV��~V�����X�yrf��D�5O��
o�Y5�
.�Q�����-k>�4I���8gɡ��bWT.�	�}t�|�,=�����'{pAE_�CӮ�t���Rn%������5w���e'm��f����bQ_�9{@V2�FϪ��:��I%ׄ��/S�Ÿ���m�#��ʰ#R��8�7l�ˁ��\Iآ�9 ��B-�ܭ�@)M6[��Y�{��e��r��c��̨�bs#p���o&��ⶇ%�wvDڡ����쪶7�2(!Ψ����\B�G3�L����1%ٮ��(j�_MSL�0��ͨ�^�sEC�\����D�(Y��$|��:J��ۛx�������[���>���-��-�b�6hG���������!S�d��4S�YA<�@��x5&%3(W7�η͐����~���ͭg����[c5u��B8��;)����^�~3�
��2	���*2e��f;�j:]�l��4����Ce��������`��?��g*�a�vM�F�����+b?�[E�z�aY����0J<C��������#0�jp\,��e��1/��;�I8�6S#^皺�T�<D��2*��d�0n)�{��L� �1�Fd�ʒ�z����q���C_�t��0�e���gSb�8��!��Z�?��(�Ϻ/���%8L�S��5f���h4�*l��/s)�ѫ@��T� �-�N�ciEp��+��,�Bw1�k�P�C�������׬�����*�����捷ު�W��+�߶�H�;�ư�[[=y��M=8$����)�b���P��}��s�Ҟ��һC3_��i�:݉	/�֞U��ֳ�pQS:�ff���w���_�Az����_�	P�� ZVpg���u���9C��z��p6T�?JjW(19woY�q(��������in�Zƻk����.GԌR�r�9����V�]��,���1�Ź�Xr)�3�E�>���KAn ���h�a� �����X����(Q,�����=?�ZI^ab}���R!`Hz�+K+��v�?��$�+8�O��j����U���L%<�!6_-�q���ᗛ�05��1�/;��/&�ej�1*��9��hC��qm(�{}�#������h��Tj��` �,~G�28�
����xYQW��C��Ǐ����\hx큽P���q#�Q��<r8z���c�|u�{�N�R�hi`�,�)�k˘�����ӟ�����h��ݗ�~��m���GF|�����[������C�|1��FVw��m���) �1���s!�tw��n?v�-�$-4���\`����'G�a�:�y����IΎ�>��/�p/:J����k�O�N��?[�$,��˓ߌ��ӌ�=��HlЩ/
n���PJ�����]M���d��;1FX���Uy�kp?RG����U�h�yAD��E)b��rH� ��Deǝ���J���3�07�����^צÄ�=~� {�nu�]i.�����8�5ix�0˰����	��I�[J��o4H���1hא�R���0ȁ*�{����@Jzg�&5��gJ��&s��'�5���a�/�Q���aD2�M-��f����*�e�@�Y������1��G��_]l�:#I��� �r�W{���̢����Q*삤�	%_�@�(�rk�.]����<��ۥ�8��\��kȅ� =0 p�:��4�f�e�jk�d;���{'�B�;
��1H[�N #eR#����!-�Wd���(h�в�@]پC!��	��!oIfG���M��,RA��YLr��I ��X��1o"+=�à6�Sݸ)	��d��	�:�vjBx,EL7NB�򯟀Iɣ����`��Jqu~�s,@ǒ�ï���2�}͋�I�B�K�2����@��}��sdj���Ug#Y������<��X��BTE��o�����\�#���	3����^���7{q��?�����<+;���0��Pp'b��3�O�9��K5�%����áӺ%�: ��Er�������w���)��(�^���%i���:�_��
��=G��VZ���� ���*~��Ԇ�Jl�0��O0����Ƴ��%�J�Yv_=n>�'1ƞ�Ǿ���Q�_8�=嶯��҃ ���0�,��Х��% �v�̡��ɹ�`�`J���N�OLn2vb=���~f<�`������|p�����⢢� �=@Y�������/"m#�޾��ӱ�+�	}Q��)O��kIs�~�%*G�A�ic�ॕ«Mj+��Wg��5�6���ڹ��1��D��ܖ��"���D=;1�޽��A�����z�"d_ͥ���"������\U��m�"��8��
ݯ1���CR]��y����)�nEQ���� �_�AbEVA�-� �l��*`�0�L�Y��,����]���H�������)/�F����cl���O�\�N�#w�r�zx��nƜ����l��W".��"_����������+IP<Lg��������ɡ̵鎿���I��k؂�R�~�#0�"s�w�f��sd���6P��|ڏ�Lb���@�ὦF�C�j{3�C]G�k�r�F��QݢK8�����Go��)�*6��I�	ń�����s�y0`��+:�E(��NU�K�Un7h*]����@f��yM��",�̾1�srLL��/���J]#���b��U� ε�ǍX���L�ܝ��CYz�T��9��2^����5} �~�м⢅���/0���ɰ=j?��A�)����7������3=#ݣxSΫSc�Y�M@��c{�ea�T{�zj�h�[	=ӫ�.% 6�H�N<UD@z��l��E���5�|@�z&\�N5%OB�q^6êz�TA{�	5t[�H����}��}�A��`�_.������s~���0jJ���m-5=wBI$�]��� �~Kʶ���/E�i̞@���X���W���9���`�����#9˂U�E
)$M���3b�T8#��k�����p����L;������c�TaEת(p&w��N<Q�p��n|�ך����g�cYx�}J� یiH�!����
����D���g��������h��2F�r;�o��GƧ�a�,�����E�`�����Q�K�(�-�<.X5O����"F�j�N猬�F�>��L@/���tb��P
��ޔH�`ya��n"�xμE�b�0)S"�'ܱ��>��+���<쀅-P��)Z��RDI�df��}B�Ul�7�W"��*M�������*�% '�Sd8YM��Q��F(��r�-��1s=9iT �7�׾��T��CV`��$���ѧý�Sr���� �/��K -q��l6+$F���<&;�B�j1X�ev��c��u|��:SM�Bz��U-IiT8CYE����F��ZM4v��(��TLgU�������E�ġ�B�M\�a	_a��䚕���lC��DZ&�P����,��y���&�c������x�j��3����K^�ݴ�,P�\��ڍ�O�P��]���MR����
�w��g>d_�?�˛g`�?�,)�U-�u�e�_E1߁��6��э�ᲒM��v��-_� 4# �@�]K�;:�67���ڧ^&���Ỉ�f�hm��#��Ŀd̷�`�=N����A�&+1e���TNX�l�9U����Be�Q�/QeݎFit��2~bx*i��R�k7r�k7>��<���ո�\h�Edjju��S��0;��{~"E��r�ݚ ��&�����y�;㹵Β/��'��7Z� bp��Ԑː�k�)���!�N���fb�`ka����Y��'��tyA��8*��V�_�u�}��0�Ǜ�b�G:~�.�S��7H5��+�o��#_pVK1��
u���Q�Β��[lk7�\ѭh���!Xv(���+ep�_!~�FL�.r�|�#��k~��\����p4I���H�@l�����{Xj��E|�m	eSL���ؗ�� k2�F���w��,��7V�t����ce�� �R[?�=[Qî��{ ���Ԥ�=���m���
c����5/�z�2N9`���Y9��.��,���X�5���*�V*m��n�,�������*�3���AG��i��a:��Xs�Ŗ��?􂄋F�o��&Ŋ�i��G@z�G��PÉ����k�U���O�jm��I�͹q��\@����VybkS"W�OZ|��|�<�}�x�h����D����i}�YX5n m
֡�Cfn�@B��,'eJ+0�&��AnW>���5�^�"�=�q<(4���m-A-��F��A�����8�Ra�r'�s�qC�b���a�K��-��*�V��:[2�N!M��r����O<�4���i�Z���'b�J��qC/>�E�9��\�T��]��cuX�v�_�s���{P[�������q��R3F>f��L��o"�Z[&A�<����d�{x��.^6�R�[Hr���^�l7Ԋu�pɄQ�4͓Qv+A�5X0�[c���	��$ϗ7��Q}d��	����N�mP*���M�b-G��Z ��Lm�����n�|��Or����G[~M��.��^�J%����2�Թ�������BD`y*��A��f��Ѽq���b�rO#��ތ��0�����_�0y��0�s�w1�k�f�Ѓ]�Ż��q���H�Qݩ��
���D+戗��V�����%�@�5�{��������Vꊜ ��f��i�ȍ܏9�)��7^�o뽏��`	ʾA�u���8ȿN��a�{`H��J�&.#�&�D�&	qк$��9j9_@�����c�����WͩnC�=�}���*�&���z�{- �f�4����D�N� �U�肨)��ĉ���� ���*gm�c]TMz���)��@ν�@{kS^K��J�+v�bo�Ȁ�>����Y�j�}�>L����r=�O*���>�'Le���,�`�z����\���!GeѢo�|V�W���Tj�vM����^86,6�����I�'h��Dq�H�<�<����y���d�c�z\���o�7$�rA��s��,�m��D�䭈8%e
�8	wF(��ů�~0�7�.Q�O2|[U[�:ڦ'�0��>�_U�)���6���4�����It�K�r���+�^.�6�Y��;I;��7��Ң\A�bLm��Gl�����Y��,T�n�N�Oދi��vt��é��?"��Z0ێy��Xm`��G�q0�h:����zl~�J���O���5[�Qy�	�B
^�
�	LNz�ɺ��I
�(!��]o�I7Ыeމ�S[h{�dX+[�왨�E$/A�#|p� Z�­u����D?�l�d��=I׍��^�����#@���ꠁ��l�c��^��ă�P�Rm�$��r��