��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����� ����m��Q�D{S���;��ie�9ߧ)������o�A�o:qlQ�����!-�k �|�ʯ�I�gr��A�PmY3t�}��`%^�"��/A@5Yϧ�a?�8��*���p�1/�XSL(����;1fKv���:�N�烋�������}
����~"�ExW�mS�p�$n���MB�X���dLqp�r¤1]��1NO��	���Ǟ�{�����A>���CFĈ���l�TI"I�Hb��Kh�]�����	��Q�����Z�[�j���֯���Mv�Lr Ot��(�R_���,š*Ld(@�v�4���#A��3��S��V3���[��Y"~{�d;(��='R�Ğ�.u�LDV����]��fok�x���琀�C,L9n
�}�q�d&�h�͝T��Ee�^�k��F6 �c?��e���FL��MȤ��iu���
3栍���m��]bM|�(.��yD@�PJv�g�D����ms'F� ,�MӰ��X��Y1� ����X֛�,A�&a=�*��u;��S������$���x�E��0�����v��70��m��H^��\kV��V�v7���i�,M�V#��w߼����g� TLY(��f�@���(���Q��D��m��;��l����B�5�z�L����w��#�����?�z�/$̲`*^�	�si@�q�3�9��y���=I��!A�*iR��Pr�R�.���:�L�͠�$SF��Q��ۯ!��F�)�?�@���80�B� )�.[�sw�"��+\�F�-�ED�4�&�J^r?j|���i�ءD��-�z[ލC�n�aj#�r��������L�����c2�.x�dηy1㢺T������5�h���F�����(6���Z��5h7� ����,k7�7��W7D�����ǏC_�ҲV����&~ں7��rB�^٤�����D���Z,���ѝ핉�$_��7?��G�����Fq�<�Ni��4�j3p�'�n�����]������4�8��ø�_=m��o���N�7�j�n����r��0��*�z�e�����C�/�4�
?C��g��T��JS���+���]�Hz�\$����s�(u,�h@b�j�HF�d^�y�C瀡������%,�����vgYz۟�`��]�p����1_x�~N9�ffB�AŸ�#SC�گ����k�.Bh~�>��\z\؁�3��`p8����ZN�w������"���WGo2�� ܻ��� ���z6�\���^��&c(���Z�BCs�$q5�%�¼s�?ij���,�Щ������ͅ��<P��brFg�JZy��8B�&��=���G@ÃV�~\�Z��}�:�F��mW��jL;
��X�ew��h�p�!R�8�{����+l�&t�O�������5&4BN�h�w�+1ʉ4d�&�aO�
/ai��0+p��`���YHN�9,<.F,�H�f������[�J�P�3o%�껦�{h�<�r��;g�"����<0l�\h��{��)�(o�|ב�����p��U�Q�*]���Jj���ӕ;d�����9���O����O�K؟��O���"�|���~��t5�6g�¡���cU��tJb��m2WJ�|��NX�\�Q6�#
Dp���1��]Ywr�y�n�J���'t��A�� �rӼ�8��&�y7��"*R�Mf8^Ȯ�����J|=<����m��DX&
��l�>�W)�|k���<*�)�HM��Z8��t�ݕD)��3��[F��T� _O�>�"L�����ْ,���̖ԁ��!I��0��q5:M��5$�BI����*Jjü`��C���%p�6�h1{�J��5X@��_虱�����A���a��YSQm�г���D���>}+{X�gD���\�`���6im�S���[�1ڢ�+�t�����T�^�����XWS����hQ�'��$�S�.�.�tNK�$DP���˕Zi���/���'h����<fD�cI|�x��]�m(����+�Ո�:(7� ����+��Yf�cS�ǣ3�i�!³����.h̶
j/}[f0ʌ� ��2v������T3�Jc Ӆݘ����6��V�*���;��_j�`n�(v/2����_��c�g���M]��GB4Fr��c��$J��Wq:��'8d��n&\=d�ȾB�u���]C��]�@%���q�N��X�%r�l-j�Yz�I�l�&|:^z,3�r	=�	w�2y��{ɕ[��L��i{��GO��8�v���>	H����~�|ȇ��q�ԇNx� �����wb@#[`�݅g�Wv�' پ"�&�ζ-)�j>n��;{��%����A;�:(m�jRE?�=9-���B�~�5h1��u/�U��Ɛ"�h�,,�#����?lզy{�XY��/���m5a��s�[�򘱉2�/u5fhH��4���C �������>��W���.J ��0�
�/k�N�@-�j���"�
w�_���)�)k�U�xK�E��Ol��'R�J�iR}��4��aJK�|O;��?�KIge��oי�g��\���s,�X�.�bX��Jإ{��aiWV9�WFKX�;�g6�"~p�����J���8&���<~����f<��	a�.8�	S���_�.���ˎr��\{d�[LxH>��^_��@����zɥ���� ��e0�\OE�(l�f�ެ�����������I	/m��/5����s��Ю�\��ByL�,�\J �k7�)l?�	����Qs)�^~/�%�cS�����>��*V�wJVD�S�8N��� ���K=�0��9_��H��-c�t��t�s��%$����~P���Up��*W�?����.�5ܳ�9�����xe��B�����G�Lto��52٠eYb@��j�)��볘{)W�����kKzB�c����j
�_����'����N���W����Zz�^�[�_��v����	�3�TmyU��-zʣ&B�E/��W�dg{�Mj̗u���0��jZw�e���ˏA�����G-a��������'�&C��β�s�oӡN�Ơhb�U.Y�s�nYml�jp�nǂ����6I��{h���4p6>��6�b��4��6�=�z�d�`SK���Q�<�2CrĐ�t�*��S,$���|����o�gG�6����]}D��� v����=���1�g�\%=�Q� `p��Ikb��[���6,A0��5��`���+w�`�0z�l��qP�cW�G�I[��.N�D 7QΊ�� ��6Z����Ee��/1�����i@Wt�#���o�H�ԃ��w&	�����+k�'|,˗8\�6�|��d4�z���Fs0�9�w�q�Iza9�CΏt���:2Z`�YxЌ@a��J5e��&B\��$�˲��M�Z��Ik���ݣ�t�C�'W�����BY��;�/�/���K�������� �ti��b�B�h��Mo�5��<ŰHC��V��C�EkY=�����U � a��ٿ��g� �VY���
�P���.���f��Wұ�)ˍ}��a19��J>~0����R*��z�o1�
"��h*Px�f��zE��FE-z�H9�p�Y�ke�g:ԁaƩc�p�c�@ ��Q2%�1
��m��M�uR>�Xsɂ��sû���\�z\���BmGZ}pMPd�y�����Oф���>���u�,��K�ܝ��
�H�c�Z1e�%����e[����&)�+�H�w���J�����}Oö2ʣ�h��F:U[G�6e黳
8� ϓ���L֮�[n^��j��z�3o۝Q$b��K� ���7��"(������Nx����/P[
t2f ��Ǧv��9$�<�����^�_��n
�>�����>6K�r�uhH�r�4�=c̖�ǹ��4�t(_.;qr��
�te$�s`�� (h<��yu�P�N��Է�'b~�;�#yၬ��jeG
��m�b�b��ɯ{V�$1���ch�ߘ�����d_Ow-l@7FC��:օ�wYU)�IN�y}G+����Myig���j���9��YA��h�e��(��K��E*7ģ�";�� D�8XX�9�#�U��)��^̓6�OӁ>s�Y�%�D����PQ_R���&
���%qn�\U�Eԏ�]��5�'�͊�$��Ǳd�S�L��i��  (f���ش2|�DƋ�9�?�!vҠĲ���PðE!�B#���4�eM�YV��,��:r�K1g����/$�e��2���7��"�ؚ�>:D2�m0|