��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_��՛	�D
������Jl]~�l�eF�l�軦��6��.�dRi
���g�h��Mw
�%tF��R���ӂ�Ӽ�z�d׃��svU�4o|����o����D� ��0�&��.X��5A����2��do���c��=��G��?��_�y��os8Q�d~���ד�˫]�isM��
yu��?*�VK����P���L\˨t��0s ڹr��}���EF��:n_�t+��Ы3h�&>�Q�7����O]�����^�Kh��喝�%���P��l�d�z�a�I�N�یy-XTtGb�-=D�D��$����D�!�$OF
�|�?!G��=��z�����^����w��=�c�
U��P|�'���D'��A�'�M�.�ǹJ6ҵ��-X6��Yd��$Ծ�gW��T�r�l9_[�}����f} �g�dK�+>��lj�J/5�6�:݅��-�x�{�K��P]�y�`�G}3�i��H��@�ʊPPM���/���[ ��
eE"���Z�ҵ#�:��1�9[-�L���(�!�i��O29��ͬtڴ�x/��3 B}�(b8��'01����������M���ڞ�F3�k�F�5\�z�*f���g��.YHk�G��\0^f�c\����क़�2 1qw�5��^����v�M��&�o�TNM
���LD���"�$�M��i�]1�&�BBW5����(�c�dKq_�h�x)�]Y�/%�Wv�,@���Dݔ^Mش<����`�RTO'GGf�r���^1�iu�*�n��t
	֋D����e�K3�")��jg��w�d
u^a������ͷ�T�E�"��Y._X��Zq�)]3Y@�����U�8�v�ܛ�a|���~S�6��V?�`���"���3�f�'��V"�p�B�<A���v|�U�x�Z#������u�ᬝO��k��_�Mnr�4>�����Yl�^��)d߆t*PC�mYI����s"�9Ż�fQ� �$ˡ؉�x��nؕ���!��y˘L(6�Ql�cu��Ȯ v���p�2��cb
�	������5/�7���ӊ�g�TXu/���4���xI�@��z���h'󸷽 �3dt�����E����dҖN=��o��}�����<4� p_�GZ�N�
h�{����#����u9f�쨆(���݀�mP��gm��87$�nR��ۢO��U
��ɾ+�PG����QҸ8J6�9�<C�\q�< ������~lK�\)Z�`!�����jg���u���yN�WP:Za8���A�P�~R��pOWۃ�3Hv]�)��3L:h�3n����<�(����y���y� S�+eO1Q�B3"b��SpM�A|�vI�����R����-�Uh��|X#}J�c�<����2���(@�=aU~��E�sRĠ���>K��=��6P\��p���vX� >����:��L��"��iw���Ky���('����! (�&�̨���ѬD�dSAh�z7�\��'[��:�{�\�XD��RsD6�hE�?;K����R�Q���I��@�wq�d�~Q+����v��T��N3в;� pYW;�����Fyސ�ȠΏm�Oo8��xM���^��T���	A��vq�(����~��EQ��-k��j�x��CA:mh�|�K=��r%Ң��&�bI,(��6�B�����3k�C���A�A����eQ�\�0F\�
�Q:uiyG�Ͱ8&��ӉM��>���� �Bc��[�~ ��qX�㳱���/��QA�l9� ���i���t����:��+��u��L����a� ��*�>����n�֓���R�]�E6~,L��;���	T��P���!.�ޟߨ�+h�� >w���Elu��EI�o} ��0���o��{�e],����oU�\�g"!�Gz��$��C�R�D��X<�ӀȻ��
��6V���~�{��a?N��&.F���b1t� ��4�0w�����qC���VC�G�G��ӕ�z�1uצ�OH.��ɟZwc$�^kMފ9��[3��y�i5����U���j1j�TZ�����Z-m&���};��(��Hᩄj ��'��"�x=�
�D�E����v���yT�\�b�����%Cs~�JA^�`,K.�;G�-�N��.z:𖲣�S�������H��#�Ͷ��Jp.�\lp�{kf�i�����񷟆^����w�uT����N{��K%A����e��劗7��D͍
51HU��лJ����?z������ڥ҂q`M�Ѓ����_Jz��sAH?��.፡l�h��9��5���>��.10S��%Pu�dB��/X�yx�^whh[!�[�C�eSޘ�v���փ���	${bS�t��Y ��e���ҝ���py����R ��Y�����2W���@��2�$;mIy�bk��y�AcN ��?��</|� 臂��>e!X�&o��\�@���
{��I�}_���_,*�o5�)n��%d*CC?b�g�[�q��o-n�޳�;?7��̶��VW����?O):�Ċ����2`����U��ݕ}�W�T�����?�Ҧ�J�b}kߞ=�H8Y7zB�mLÌM����e�=l��-��X�o"�	#��h&��gt�2w��]��Ĳ��f���?-.��|fȡ9Q7Ѝ�J�4��Ih�o}��/,68��h��d���W�X��/��'�G,8��L�h�&ɲ��*R:����R%*(�=�T~�� ����di�������O�&.}2�a��}���x<c��;�-�z#��(��`�/l�V'��2����0�5<��Vq�Z�%��Yk���^1�_ԢI0����^%0S����-��Zf,�4g6�6F>�Ȼ���OB���L�*�B�K�Mȍ��3�x��k���tDT(�f-h_��U�Coݔ7H۫]�
nP��Q�MP�Rb9M&��i '��	�`�G�m(?���I��m?as��� &�пo� �yq�Ѐ"�t�5��{��̖�ԃ�����/�Y+��E�U*^���E�Λ��Y?k���g����
}	ֺe�(<��=�ASy~ђI�	�/L^C ��]�]!��n� w�鯆�9�hQ�&>K�W����9mU���0�M�ik�
��{\St��0���_E&s���)C��N6�0�ҽ�P�����Y��y��/����1��$9r�I�(�X��(fL�ȫ-�G����A��f�\|Xm�xД���F�S�2�����G��r{5��u�ۼ���������("�-7����X��%YĚ!Y����HS7Ja<����~l���a���J�9���k+���Diw�ԙ�����(�a�:i�_�Aǎ�%_�e�edZ�%�7���=z��?�����1r��̈�I��;�ލ����j@�qU9:h�@G�7:޳�1�L�L�G;b:�A'UD��5e!���ka������$Rl��>�2
i��JHJ[��R�������u��U"�+��V�V���%4��<�٘�(��0���p��&~��;qd3.��C����"�b>	yY��E�h�F��NT����ے��
T����ع�	��FJv_�?iQ3���s#����=F���/+mc�w��>k;�A�ܣ��Q�Sk�4P�]��B=��tZmLw�����l�`�����{�i�Ca�3�}���&z=�Rm+{��J8^9P�vL�h�V�YI�cL�sq��D��T���0�2�̂�0)�(�7�T��O�rV�s�� UQ(�~뻚g�ŨV��H��E�9��f�����_��vg��5qV}��	�Ǻ��-��޷��v]`Id�5[�#ͩ�S[ɕJ�J���JhQ�	��!|N���l�x���l��^OH�r����/��
eu %:[��R�%+.�2s��nS����(%������S�A[nI'�D�'�w��$��Re�Y�K_��nT��wR�t��uO�ְ��"�
%���8l�[ �2�|~�r�h�G9l�9�n'q>,l�K%?���5���iZU����,G�&\��tQ�o�QD@���IL��t��$7��U ��I%�۬$>!s�����lmh���v\PcXҮk��V�I�|���� �n�KeU�C�XS=a�A;��-�ٝ���q�$��yA�|�����ޚ�0���)�'��B�k�W��^�V�+��'�4t�	�?�R���>�=�q���~;rW��L;��S����ה�5"Fl>��9�N�n��);�S�E���\��)�%�o!)�VkA�%q�L�W����
w�	�0_��C3pH/%���f6���<�p@���JHt�(3g������4���6���k5� �Q���C4��@��P�X�h?]�00�8!���f�#��ob�M��b;����D1Jj;�&�T'XEZn���)��3"�D��{a��0�ʗdQU��ob갊Ze�Jw��o�F���� |iڎ���Z�"�^��+')D��v�ē�?���2�c�BA�{� �c�^�ȁ�oHjÝ:�� I.���5��8tN��_|�`�;鸢���'�	)��Á��r�Ax6c�Zqf�����nu�7�ῤ����Y����Z��D�>+S��]�op����
�d���t�Q�;?�%=�0����q�m�_ 
x��#uI�GC�Ϲ��I�~:�@�X��T� �GES��$����-�^Y&�b9/��)�J	��
�*�{5�|�;���]�������`���~x`���+4���*eB�OwV�.J�3a���j� �LaΊj����}��e �Ie�!+8��Ex[��ѼBW���K� r�������C���X~�,��Q���m�0����FS��}���$��Nݺ�,�׭�~��9b�8n�$!ε�-P��޴b����8��q�Ӂ�_�S1��ű�or#���b�eu�2#��	s4����.JԹ�Ӗ�i�dU��?Y�QeTr��w�C���2!$09(�c�c��-/�Հ�w@��椡/L=��#11��1����2�����`*힖���J���$�ߖ^<sA��oF�A�W���7W�"T�*��a[�����Xo[���z��Ga���ɥ���§n*�?%�T#�~��]�^^-q��;�n�ˎ,K�נ196ŀYU�U�����TJ��h����:],&�z��x��f�(�y�Om�wژ�����=��H��`�N"�Q����\�,ԱU4�4%`m(�.3��U���~����eS 㼔����\mt�Є`���.#�G�n�뺁��u�1h1M�d�����3��x7ý�3VT��[��7l%��Oo�CГ/ڭ]����?Hp�s��u�.Z���p�{k�7s��"�g��"�񻘱�M��Bm�L,��` �Hq��g�6���T�Mi|i�J�%~��ȸ���k��E�����+͆���l������iG7e�I�-1[�mߌy۝�)���(LڭE�`s_z��IÍמ��o�[3��~��y>�*n^u��9x�~��4ƃ[#Ȫ���a��,����=F��©LZ�)���,T�Q��T�ө�ߐ�]��t�JfqK8I�M֯��W�/cIs�'0g�&�?��E<*p<}�M����a�?�}��#��}z��G�@{z���`�`��੐<W�S�
r�a��W��9����-��`"�j� �EH����a^U,�G�
���6�4�U���˃�<���p����+�䵧=@p�'J�qT|��{/��g"�/�*h�Y��`���^c܇*w�E���pr^�[O�"h�J?�^�1�����t�������%-9)�˛x�+���Lq����4��y6U
�%��Z����ˣN��n�QP7Dx;�ץ/��VmY-+�ѶK��㘿��`���Ry�y1KS����Y�9
L_�����4]�/CD��'RI1
+گ�n D�����0���ƙ��:8��Ǉ���)��m
�ޒ��_sM��Xnb�7HI�	��&��$t�8ؿ� ���ѭmG`l�}^z���/��ҹ�x�f�
�
q�7�6n�����j�54�db��?����/�_�\�׺�����;d?-{Kx���l��1����C�wC1����yG��ռ
�1�~�^��r.��\�鐍 ���.Q��g����h���h�O~.�d_H�)��24�J$	�-][xb�*:\Jg����Ҿ�l�� �}"��t���pv��Fe���4���>b��B�o.�&v���)�� G%j����D`Ǉ�5�,**������ɓ��̡�;��h��{-���r&�!�op|"@�n�d'�v>�ʠ�r�z6@l?�<y��P�Vs$�s�<�¸�a�x��("�p�p������M�D:�r�uyQ8x��4���-~��sQ�Nl�۬UB��v����g��� i����H���
�!-���P��k�&I#���g1�C�>�a�a%s���.(�!=���m��;�M�UW�Q�~:d:pk�-�F��*r瑦/x'����	�´l>�o(�I�$�^9N&6�_�9���ʓ~�3d��($�"����4��7��Q��a����72��R%��&=,�w�&�d]��W��4�Q{�[++�!���j��lxy>3�~��T���E����,:i�G�D�9�<�Y��<��Ch���WV�B�"���z�Yj��H�W2��pSj�X4C!�A�O=U��W���~,	���MG�U�����:[-�=�k�]�@�L��k��#����b��;����T�������%B�xk|D�;NP~��~�>_������#Rx��@=/����L�Z�W�=oe�x����l>Y=��`K8%lA`���(ZG�} ���чkLم��0^�*��bq����˕�Vfa$t!J���w���̄�_���b�r�V�,�/'�*ˬHa��$$W6�T4Y�ي�#�h�����#����"4��1���y�e�Ā�^RA��� W&��M�������?H��B�כG��>6��E�z5���I�s9\�}�>������ِX$EJYNf�ts�_��u�
��a;3\�(w0��iP�$O�c�G2���DD�)�R�7�3���K�ԡ	p?_��F|`����&o�{>�ˇ׫R�1s���\@f-2