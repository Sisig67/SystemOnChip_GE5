��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��E�a� �f�9�?�p(�����L��R�U���vh�����O��כ����U��\`q�"���������v�T�Ԃ@%kpZ�b� 
����D� h��L��`f2�M�bIْ�Y~�A�֘V�#;,/�@\��F����`��Ԩ0G@` �{r@�\O���K�Ky��-��0��>����`�F�����9F���d�����Cш[�c��f���ĵ��ji)/����� IV��N̹���.~~�/FR�ӑ)��p�K�ħ'�
xGS�})��!ö��I|BP�Io����N�@�79��Z"Ę0yΏ�+��-E���"ﴭ[�F�-bңW�hoNLb5��m��"�s?���-�4v�6�׾���!��1���"�W4�`aBy6�R�张>uD���T�tb(Y����:��<�N� %,�ꍬ�m�0d^hRY�� ^�z�lֳ�`
k�*@Fh	 P6�i���<Ӕp����f�m��v�)A��Y��w��jF�6�c{%P6)X}xl��P$�`ݢ�S�O�"��7��E��M.ɟ�� ��OQ^�i�j�.��ʻ��ѕQm�5
���iI����*lXp$0G�khJ Q��/�e<��@�FKK��'� �g��"t�>�δ�X�A���F�.�Vt��m\]����w(�D�@�W� �J�W�2W<#�&�q�\%��ν�γ��o�_�T�P��",נ�a��דg����v�����ڻ���d���J��
)@o3ϾV��V��]�8�w� y.;��0XƧ�sc7��� L"H���mJ��TA$�	���Q��n�E$uF�4�UJ������g� �go������ƍQJ�u���ʹ��E�{�=w-`	�j�瓕d��DWD��>�B��e��Uc�Z�*�ԅg�0/�])��1��c��C	$���\�Ri�؇�.�ioz<�6��'�L�1Va�G"���:d����>O,���1ɾ	�y�ڛ����k��H�#Pe��Q1ׯ�2a�EM��i�7j9X�����Ƒ'���mq�gՒ�}Y4�coS��υ�Ȃ~�H�u�^*D��=Ď�{F�܍���^��!Z�g6y�~c<~�%�P*���Ф����AV������H�Y,��n���[#���5�����1,)?��&���P�ފ����N��z��L�	-k��xÆ�s&��MSa/d`��Wg�m��ȅJ���j|t�z�;t3�Fl�t�������������7��idi�/�����Oۘ�Q�L�WV�!8-!�P����xx�5+^jPC�8�óHGuV]&{~��Q��1Z���j�@��I�븑Y��! �x�A�{r5�e�
}�-��P@�U�ȳ�ɓ��~���UZd/��l�,.�'+|�(���b�}���Z2~*�;��-1��2�ThG�t��Py���g�� ��Mc��v�	�%Sb)I�����R���ۈ��i����%�Q��ng(����`�{�ѓPD)����p��j���`�:~0]�:cߔ\�+X�Vq�V ��R��)�P!��D�mĖ6n��'~ɏ%�.�y����.�&���uy7�� 7@��W�-���O�
HX@X5<JZ˻�.t~��K)�ui�[�O��
�����^�j>�58������e뺝��F

�p��ﭠM�u�����U.Zkf�MDz���3]��%E����*q׹o�Z�[͢���a�)ij�yA�5�8U3'������#f�1��Qo��9�TDᱶ��uoG�1_-�7�������^ix�ܤ�|����mQ"X��3�{�7+���:A�D.f��ʤҟ4��p�*iTS5��KRq5A�v0�6M{�EJ��M�\KI&��ŅCu�)Ydh/��6�{=�+������I�̇7ـ�����+&�HyC��v=�D�h5��2tL���3GʎU���J8��z��Xa��ĉ�p5+6��\�0��ܝ���k����5�|�����i(��128�$\>�N�-.P��"೷@�-��>.�ePj��B&Gb�kɱ�o��@��l���&���������jYx�t�6�.��YR�yzN��	��W?!Wp��o��N�����`���Lxo��;��O�.��?o��"�������W�{��m�
RKd�U�D�V��/�w�S�)5�N*Ċ�X%�SQ�L��CeBDI;ծPf֏���k)|��H�,� �7`�J�쳦ı��U y4�׷󙢓rf��G����<R�y%��������Q��],�b���"���@0��C��Q��V��뾸�d�Qr�i������=�*�$������&m���?����ޯ;!Ւ���Πn���D3�@;�ԧ3����Nܘ�(�����Ĥi��R�-ᕓp5e�hK�Pk����"�Ϯ�Be#cXX�Wp���`(��ƃ� 促F�Zr��'F+��08�ނHN� �
�]��D��eg	���&bH+���ZDa7]q�\��*�y��sax2�����Ib�([X��t���������/��j��Z�rˤL7gŽ���R{�MO��%�G��|y"��@�Q�O��[�2�Ϛ'54C�l�W +9��Q�-��[-&���a������d��'*��b�l�Z姂�Z�d�v���L��N���K�=R�rc�?�E�w�����/�LN�e4�c�p�A�E��s�MZq��2����Tw�J�&/�̚�c����*	���(����z��
�u�p��$p��	�s��:g�Y��t(��U.0"���,�L`=r����]41Um�gԊ
vӿ>�7V�cS�h��E�ۙ��*�<H[��a���d�#Q�8���G0mx �cctrh����	�mBq;���;��]������n3�Yh���] �Ĩ�,����#�@��ϰ�qG�<�y.]�h��Ja�@c]�כ!5k�R<ԴY׊Jl�7Gv�WGo�H;�����yi�j�>_k'1ӱs�Qq�)�a�VL��u�5p��|�}�����n�Um���%�sx��C�7bl6�A�VP�Cm[2�����x�W�����@j����A��-����Ѿ)�k��5�6棡�����.��r����������*��L�:��:�u��Gt`6�����!��E�]aN�R��UʖA�ޒ���n@���,L����d����	� �����#:��.
���*�)�xCJ)���R�#&k4⹅�--M�
!�1J�Wr)b�����"�96}zU��ZuoY�ї�ڞ��\RPU��w���2 b}詧&~������Q�1Sm��i��p\� Jw��J{kC|i��iqI���:'�ʴCXKg!xV�JLё�VD�N��1hk���I�>�)]��Q R����Sc�8���`��3�0��V���"@�G���77��|���.p��=$�<yB��$�N��9D���{��ʲ;��>��TvG�8���	�S�8��A���ʖ,�F����U5zAK)s�~OIF��׃��+9y�H�A��>�F#�6�⩳�:��������;DLe<{��%�� ����ƕm���ͼx��}�|s�le*B8��	��/3�
����M�opIł
y�����=ti�;�b��I���FR�*u�|��.*�n��B3��a� (��(~�4�)�օ�O��f@�J���1��G�ۺ�y��['�5��?�!u����K/L�*�.���$��K*�9���?�r@Яpu��Y�����PH�^i�� -�v넻�U.H� 
!j���+���-0o���s��m�X%b��;��u_wcgk��%��7��I�^�ɟ���W��X>f��FAj�o�d�����A�AY#%�����Y:m��2�W�H��2���"�h8�*��W(zo������`@M�������!�bkgf��L�I��IƧM�]<B�:�%'B<g�y�����]\^|.f�  G-�%����ڬ2����lD !E��a��z�k_��J�*�Mʱ��ʁ����i�ڋ|!���X>�^�"�{� $ԇdM�? ���u��R|/��ƔMе9���F��Ϝ���y�`�Bmj�1�y�+�O9��ț�`��o_�V����,�����!�2�7��5�U�!�<�ܕeج��⥉r���K^V��	@�����b?�	�B�U�-4I�09���X=�e:�5��e��	���k�%�6�Qa�x�1l�.6��`wd�ղ V��M�]�S���p�\��(8K�V/�-+˥����t�UTqf���8�P���>9U��ibReE��2�J�8���;��g<��M� R�#�jr��ƕ�I�d�d��� �-��l[�,;��`Q���U�?�(��YS��i�"ѳq�1K\��|v�P}���X	�w��1�
�;�ޏ��5d�1ae��ސ��{�T� W�g
����6>z�kr� �	a��fɻ'ѹ�������sg^�󆡟pA].g�,�\�»��,�M5z2ȑ�V3�d�]�������@;��b���=0��K���F:��}�>@r�2K�k)��̭���v�uch��=��IV�S�E�7c�\ �g�zf�t��=���Pb3-8T7%��]�o+p�łˑ=�4�3�1����ֳ"�& ����1#��U�}���q�׾�*`����������g��vގ=��m�!I7g�"LsUr���kT!ǝ�v��9ޚ3�`kj��,�TQy$��u!8�`�Y�y�.S��t2� ��~zw�N�P'��|,v�NoW�qm���w�(ch��:Jz�J�u��_��:�S����Y��̗Q�
|w3�����o�"����w�