��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�djB�D����)gХAIL���b�)E�
�Љ��띠���H��la��2t���,��u/j^��С�0�������aO
0+�죪�Tһ���RT�8�h��oZ�׉e��� I�X?F�Y+H��[q�����Qݠ+Ξo�L�%Ô�"�z����XHb9do"Q��|T8��T'��jr�+\�x7<�`�d�7[�������v�A�ؘ�Ђ��9=Y�?RxZ�Ѥ�^Q���J�E]��j�ꚮHcN�/�'[h��}z#�*g�I��:tl�w��^,� Y1�/R�I���/m��ǫ�	���N�F�8+�V.�I��

PQ1)������N�ۅ���8�ߡ�uk���:k<������(����}��n�QB��@��1�|��~x��CT�q�P* ��Q����I1`g�A��TEO� ��^�(K#e�X�U4P���Q�Gߴ�٦��ipɁ�<5��'-���3	���˦B`�i�Uh�"��ߜ�V5����ya�8X��	3XX��)c@3Ӆ@f� J݂� ��͕D!7JP���S׿�$����b���_�0�C��	�������׀�Lxbm̯<,]F�/�	�ZN�)/����T%ս�*� �ix�ٰ�St��ɜ\��p����^�M��,���5�oG8��'o�e����,v�����9�b��b�_�2K�^���. ~��mJ�n?9D�=�&A��G�\c�]up�Gs�q�'M�>�|_T*�ۃ�ߪB]6Q8��^�m~��4�0lL�ˢ�%73�M���Pk���E;$��;S �����5M�4}	�(ȩ��;qtH�и хH��#$U]�nYF��q����$�_f��n���ٕ�c_�.��d*�
d>X�,H�E���Y>t������7m�S�r���o���z|M�ه��	9��+�@������YXo�ݿ��yV���,uc�8{�� ]m�A4�v�qa=��I22ZM�0�߭��"~��I��a �YZ�g�w��s�>�d�j�N�M�-�f�}�x_����B��ɍJ���іQs���̹�C0�xϢ��C]ԦNvU�8ք'��æo2^�,W��@�� x���1��e���a�@"���:��=_{��˲�?��;��Ӓ+Q��ii�'�tUm���Bb�����u5s]�ˀ~&P����S�m�/�/`^��"���2a�Ԗ��t�?g.�e1���JM|P|W"���~ӳo��k��;Fa# �~��KQVV�6�E�~t����P�4�	�Ì��:5�	o0�t�Q}�-���pgE좈0<�m�$���WJ���WY]���S�4.u ]o�x{j>���>�$����YZ{:�a�8=��j��C#�b�{R��h�1��4��أ(fn����2�a���H�JR�5�ELE���,�dR�� [+}�E�S���W���.oJ�@v`��w��y�:@��:�O�x+�����fm�Z�ѿ�Z��a#��4��Kɖr
�:�H���	�������9J�\/Sdh�٧�e�?����t䰈�?����
gL�ļ��nU��9�j'%:)���Y\ ��X���g�-y��%"���;�';ӧb�BS.���~P����|0k)&sMֻ��A�j��q�<�={�����z���Hp@A�-�e1:X�������I�B^_�	�0���A[]l�_��Ji�i�d(�X��e����ߤ3N�W�xϫi��	e�[>�����!� �69=���&F#tטּ_p�
׋"�&�8�?�w�b@�k&�(-5���|�q�� :1�MK�s��:t�PCY��L^�v�z�1�.���=2D`Nuf�%w9�ע���eDJ(���`.���z���L؁��#^P�]I�r�>�1���-5ܣ������Q:��@X{�1�m�U'��8���|�%���n_Ù�]�d|�e5sZu�:M(<���ݕ�����4w|�����O�Y<��)�Ch�f4�~M��@�剤 IBF	Պ!~@_+�B'�A1�=�1����5ȸ�^�4��ƶ.�Ye�l�%�d���I��(�}y���7�L'͙)]q�{��C1ԃ��\#Ɂ*>���%�Jp������i�-��'n���j�w�.gf��V>WOk���,%���e%pp����5b()�&ݽ���?-�7-#;��k���R����=� a�A��N�צ ��y��ɶ�TStH�1>g�'�Ԏ�y�L%� �{Ӝ��R��Ņ<t��t-�Fq	Փ�oz���J$�<;����n�]�k�:�2��;}m:����`���d�/'�'t���ሓǔ�L���P���| F�*�^:p%�/9�4ӰW�0�����	&ֹNB;��߬���ᕣ�A��u@��R��^|�<'iN0z�����/o95[��mE��"��"<�4^����U��<�����#��(��`�1����D.�|=�6L����G�#s�	}��x�6�6��2���쑱�aO�*����며(]�{C�&�z�6�e�\u�ѲO;��d���1O�����LY�N��#.���YHt�}	�R\�>;�)�#if��9�u��m����@�Q�[�f�5��I��A����9���۩O!�gs,�f���Y��3�=��NM8E�Z����(��Q�'��m|m�oo�C�9�Y�jX`+m̢���?�\��� ��:��1��l�$ uh���%��M��nO�$X4?�x}�3+c��3N�{�NkG���&=d8Ny[`K!\�	g��U��'[^��Rο�Xf����zS���N��ϰ�w_x���\�����Nn ��^,?� �D�I�ߋ;6��` ����h�� f����J���׳��t��*g����G�6a�[��[�n����C�/��ry���~D|�S0)��O�8�\����J�s�I�V;��a�9�V�J<��8��������lX�gKy�Q=x���e�n�0�\f�8_V�;�s��}����t�<8�<ף�0|�V��� �|�w�Di�+f�b��A$�L����?_�{Z�6s2%���'I�����ݺ��7�Ӹ/	��h���x����,���O�cv�G��WgN���k�~z�����6�����E����2������f1 ]���L�F��8���1I�Bq+��4G��� ��O9{#D'�o:|����sP�X����wD �?�>�W�	e0���O��^z���n�`
��Rf���#�1=� >ԧU����FŲc�P����'}��;F9��;潚=3^�: 4]��O���<���T<nR��[��-�h���Π����V�}�
�������	o��7+ >N&[D��$}��U��+4⑳��gج���u�$	Y�{e��"�x���z�ٵ �$�"�����"��|�fР@-�n��&V�&o������1"�i���"d�<dH�����W[$W�b"<�Y�w�{�*[谰��A�W8�Rn�j��]g��g6�������������[�U�S.��4(�4�į^�$3�}��|r��Ϡ���"<�_���l�9\�A�-1�l3Q%�G˔Τ���j��M���ah�܋�,1D�!M�6��}�^�q��y��� �d�s�r��iɿ�u�|ɑ>�y�͝��O��Q�� ��::�����&(�~N2Ӗ� l	��#
=�d r���q�#���D|J� }]�=�pgؕ�b7��5ဟ�/3�mdbIj��%pq�Zw r��{�>��4�M,.-#]��;7���&�k�,�̔*�d����o؃�@�	��eD[�6%�=�w�7B�{
qc�sD�����1�n׶�o��-��uJ|�#H�:1��[췌�C<MPh(P2l�}�HA���p�|:��͓�K��[�oMKFᤞL�?:�
\Nn�0K���b���j�=0\T�CYf*��#�\��Is啒oLOѾ�R�?��yLNt]:d��;~��Z#)��T@<9P�MN���C$Xyѱ �}d��	�Qn��z�p��T|�VP^#�i�	Tc��+'�/AϧYFAS����61�9�&���qۏ���(yp�� +J�q�	�^΂�%
�5��Ì���nYG	G�,�99-A^�c�~�>��:����Qs{i���~��S�2�����3Z[��0UG�ˍ|3`� ��f��A�!���\� @
2����!�S�K/�3H ������ya��@3��d�n�����IѦ��|�&�rd����fA{�4f`�t�\��E��_'::?Y��[���hm��ާqd��^ήJ�˥�s�zN������T5cn�C٠�.���jc~lv���k'��)q��R�e-y�����e������J�{�^��:2X���t���j��)�_�o�S�������ꊯI TfK �K�K*���1	���5f@%�UܭNu��� `��&x'2��L<�� G�8=/�Thk���J�_�/��ÑD�}Q���/Ƀ��6������|��c�$w|�s��r"�/���y� ,�s��0�s���j���U8�Ť�/�=��+k��o0/!6٩a�0�钂n�*�p+"����l���N�״(��Z{��6/r/`�>u�<W�@]e4:٘�� �7���m�h��~uQ��!��飳M'�G�R��4�4"����R�  �S����!>�{"N$�v��	�Ǽ5�f�f���|��"�QO9�x��5�י���Hz?���+!C��������!5��~$<�p@lNa$��X&��?w2����8M>o�n	��*pu�s$��-�t����N����=Q��ȣ�Z�j�F�H�n��Y��������}󣡂��F���/�'�\����m^���QMc���`+�8�5T��x��I�>�2TI'?�jb�&?�S2�9������E������Wˤ�nւ��?�XzoE_�<T0���'݂h��ȸ%[��ky��k��w�s�b 9L�[X-Q� [�v��Q��?	f���SA��mvl��TXU�o~LR�;��0Q�����2	MǑNy�Pj>ɩ��RY�lВ���5�7���Z��?��B�ٿ�\������e��g~�B�פ	�\8U�k��i�1��WPQ�h��jC@�@N=.��A�d*z8�������
.�iS q����9�T�0�W0fqD;#�;_�$��nɂ�x堍��zw���	5�� ���Z=-�R��`���Z��Э�u�SK��]b����e.�֣K&FE��K���u-6��#A���O��\�/��}��$�̋7=�����W!꩹
���X{u���D�``g22�0�\_��<c>���`�v�Xm�AS���*/��S6Q2!����<)����ry�K���=�^�Ӝ��hn|�V�V>
��͝ք$��1C�B�"t�����\�p��٩*�B�ݨ��������h�# ��-�Fg�i��x���2���I�����ӷ�7�3�Ws-���[�|���W�%����Q�:��JW_ʣ/�_�C�>,�*i9�)����ӛ�:
��D�z\����>xKy�%ds�h�ݙ<�����W?J'-����r�v�ހ�A?uE4����C ?��2�u|�	�m�On>[(��.?���
�m�3x��a�l8O�<�v-��&���8��U�t0C�/1��mje�L8�0s�7޼V|�bKP޳�qt�.��w�HK1�C�����2�t�,�hVȚOpFf��ɺ 5e�L�Y�#�A��
/��e�|�(V8�z�=
��b��Kr����y���)�ɋ�ch��gP`/ץ�\;���+~y��;�
��f_����X����d�Z\��Ǻ���|ց�e��P�y[
�<\ܙ/Ia���F5zXhI����ӯ��`GRl���	���I@����7ځ��&)��>���Cǂ�+�(,��ƈ(J��\��g�Y֜�#Dz�}&��fw;t�(@q�����a�q�XS�瘆�ۙcln�.[Zҕ�l0Dh�p�!�h�Z�j�a�4��ҿށ?0�8���o��},�/�|�b�\�a���!�  �|V�zQX�z����	�9,k���z2r�2�o�W�`<��2e�rM���<KKx:KR]s��q;�S�z-��z��F��"���
�A�;���)�|4~����_�C�h��,yy�'[8��'����#�8���㘝��A���+xy�L�7UΘ�A�\B�٣�K1Z����4���Rv�� �p�c�3p�u��G뼤 ���΁��"�:�֮yO���7��s���l�a��D�c/�9m8&��	o�t>�}մr�i�1n�5g�[�b	s(]9��0
�ϋ�LῗHmE�qg��5�!�cT19-�����7Ќn%����x�B�!i�i�7�ѫG(�/Uy�f��5���r�β�45�����4�� N����������W���K�ߢ�a:l�Q�ݻ�D�>x���+�����D~l�ݬ�+�Z���L��Cr��ӋE�$+��9P�r�b�~�,b,{����� ��';Q����v\��n��*~As���@�s����,����p��[��+�-f
���-4�Zz|͟'m2�e�)٩[��@�AQ%�Y�h[x|��_-���-�V������%8��X�ާ���i*Q8s���`�<q:BJ��>0AlE��c�����N܊@-����ܡj<�F!@~�r-[X::!��d[JF~d8�����z�/�}�^�E	�_k�`�������50��i�7rw��T+�Z3ԚT f�����X���{�Ou��||�bcYi��J�?�t��+Q�o}Gg���FC�|��䱄��	k�C<4�epU@���GwcR�@rNR����|�$dԡK��D�#��h3|D�CT���	���<z�y��b���D��C�7�b���A�?��	�3�^�عi�� gV
ج@*�l�B�k��k�c��j�x"����f)�pv��#����vFm���궮;��'�L�s@���P�ǒ�PwM�*���?��Otb�Cx����LUS��3˪��
�!�	���Տ͟�����e�'�:l��������̵yos��8t/�!j@ϜJ���#5��PW2�__��#�\�-!ɜ�v�?�$���Y�PvUU֬����$ln����8�}h ���I����y~:�KfZ��q�"���B�7ϔ�h���?��X*�hQ��ڊU,N��M�s������cJ)a�X�4�)=���wn��`B�=̥z߈�����J�},P�$1�eh̖��hW�713�g����5;|�/�[H�����3��\���y���ȱ��<#�<�R����楶s���)�hd�BE<�>�h4�e�?[�\���g�H�*�B����A�L�#P8�2��e@-Nr���ƈ�'4G�z\��N녻�T=
߷u��w�L�a�t���)����e���u�W����)1M���܊'m�p�^E��.�ǜrP��~%S�v�0�<�T����1(�No�[��2x�[��7�`�(�6��cU��P�eĤ���<-��2Cjl�}����{�p�P~1m���Q��M21$�0`�T�pn����y>���!R�#� ��f���n#��V�4�� �)�e7�Q ��w9L�ʧ��/��SLsoK�G��a���Zo%o<,�FhU���-�^��|�E�:��I0�f+D��\���*C��@NN��.#���׷9���ށ���¯�5e�!�J����HA3B#��m �O��/�ʞ���6:l��!�в�l�,�)�kf�DN��`c�]���u�[6z�ڍ���.C"�¹w�_o�.��e�Mp��Q����SQ�Wp���S�X�Mg���j1��7H�8���(6�i"a^[F��	B�H�i��~��C/��C��zHV���"6����?�����53�"�s�I��Q}h���S���Uc�)!ʋ��ܹ�~�I��^f�[ n�L�<Ԃav2�rg�k��SF�^�� H���x�G�E({6/.ޡ�W��Z��;�q`�D�2�}��!<��$�xJ�ߡ�m<�1�G��O��L=���	��e�"AS_�T���U��ZS�e����s+���?u�����Zu�乚9�q�*Gf����7]�Cv��W�P�;��db��	S�cw�������u���D�j6|�۸Rb���ʗڀ�r�����:��	��Ӂ��;���Ӝ�G�@_1�B��'~��=�M��l�+�{��}oBk�&�8*�U�u�f��7H��µ�8��Y�k����	�R���W,��b
���_�j�;%(a���8��2�M�{�uT�8v[�Ǎ�0R�|���@�2���$�%����Uq��e��<�Ŕ��n�Q�	W�4<����A(o_|�&o�!��+cq�@apٸH ��ę�IO�����O��������tc�	��܃�g���	lDw��+'��'��Hr�H/�A��C�s�1�4�j޼'�m�#�uzn�}t|����8��E��Y>�h��S>�.���e��s�9���� ������(�[���/d��x�[}�Z���^�qu�yG�!��qGr�WK\p�����=��Τ١2�F�{�����D��)q�:`�FJ\ֳ_��&���Ƨ*�*vu&��PA�J�g$,��$+�fA�*�� ��\�;P����<�!�}���mB6y|z.�t��A4�P��L�q@��s�(�9�M�T�d��IKnf�חMP�Yz�@P�}_��%_#+d��L�]�亅�؊�O�Ix��@r>���-l��7�=�2gD��n�2c��H*�f%�.Їw�I� D�Oad@��ԥ�	�R�$`Vbj0z��ݨ�T�Az����G"�K�*Rom҆�>�lj�g�5�����
U�`�Z@����Z>��xՀܼ7�4��&�͒ ��8m/�i\�G}�#�엥yJb�"�Ł����Ԫ�W6`������޼���޼��)g������Rj����[+�۵�*�x�v.�����e]��W6d�OM0��X�9����/��M�=��io��:V�����@���M�.a��y˖@�$dn)*~?��_�Х>(�'��g��>ɬ��E�$���MV���C=��H�B���H��8ۘ�5�`3�fJ�=;���I�W��J�!��D��j�殌���,��b�V�@d�^�.�������<�A��ኀ��L+	*@����4���!�\x�Q�ї�(�����&R�C����2��VqlO]�t�A����X���v_4�%Z*�} ,p��U��MT��ö�m�gJ�6���<�H��g���?3ͼ�4b��������|ؙ�b��;��>x�.k��-H	R[^�Ph�oo��P9���I��(�B1�k~����N@�����p<�פ�&	M��%�����eL�&� �v�+�GfXm���ƪ+jS�8묢�_'��������|���ûK:qT��+����g�	D�A�0�M��!�]�e^���aG�� ��ܐT��}|2�L� ��˓��@c�2��熜�^Cw [ ��JK��}d(��LC�Fek�ުe� ��לcX)�\��ub��S���:.��"+qH����ob�P��"��$j`�g�}c�(ID򻿈���yFS���)��
�d��?$�`���֚:����g+�s��7��3cR��^Ч�V���6�aa�܍���x)e�t��Yz���СL���0�N2�N�����ʰ��י�9�h(�{����V�T>�C$�*���?�M���癅eQvy6��"�����N.+�fsO	�4�AV���]@�z���w�e푊�l�sm�ʃ?w����~w�������� ����X2�ܲ$�Y��%ғI|�H/�ݦ	�����\�LUB��{��DC�� ���'�B�m����T��$N)��� ^�u�;8a��l?����wƍ��O~E#���6�ݯ9��Y��)����9�'�4ޢ/�����7rI�_������N�c�z�bMÊ1��&�y�y���y��cL[��]*րyHI�;|z�-FE���	@T�Q�H�dh�����W���t� ���'����zpo�d�M}�#=�ʴ�����{��lz/������r��!z=�"����ҘKѳ��vjw�-�5�)�T�?c� �&6e.�p��Y�!k�RTs��?�c�E�#ڎHQK��I	/����, X���d��gh�e��пڞ�\�m3�m�ǠnG�Z��������z�۴|��Df��s94��L�X�VZ�Ő��|����jK���'�cѳM�q.xS��϶S@��v,��\|C�1O�o����q�\���� T����/.x�B�Q(nǭ(���DL!�B��m��F4�������|��5�s�����(�q%��~cQ�d��&��:�*��:�@���n����`M�2s�Ɯ�|V���1ޚ�;������ςeD]�u/�B��/hsy�愇��
���
 ���\F�^Pd� S�)7��[�����0� �����X���2�1r�S�N�:Ǻ���d<,yZ���"A�$�.�g{����b�0�zb�����{���)�{,AN��ݘy�Z�н8?���`��Ӯ ���z�T�鏓����en�\3�d���oP�G8��R��7�H:�8�Ki��<d�րT�cҽXs��3-Sx��$�'�/|Pg�JE,��#6�mda���'ow�F|Ξ���J��.5��{�����mT���l�XŌ�%ty��uz0��%�A����iVT�ݍsE~A�����7�����a�DR�ۋc�
�o��,w�؊#)mBgܞ����ynf����z+�7D��A�u���5K�_ӥ���_=�|'��9�G)[�����y��P�ԉ��Ka�e {�����[F�+�g�eMK(a�K�K�y%��RA�]�/(���ـ�^�j�𣏁-3�m��l������S	6Y�T��_J[S�L�1�� ��a}���eɐ	����w��sn�k}�(�D���֍����VG ]?��͹�����}���]W�A;�������X�U�	�|�6�.��E(��X.���PIy�QX� ��C�,L�
�x^y�-�Z�A�V����^�W�RXDX��b�nrY&]}�r�d�0�굊�{���I~#���d}&�j΀]�NwܓЩ����N�}����ɋB�?I�����+��N�9Sܛpv���u�Do���p\ƻ���ޞ���ez6�̨��QN���;n�(6�<�7'e�uv��܀��E#�2��6e�C�d���ö5.���(|I>��##����'�mP>f��'`��!�/Z~�I��&A�ĪMn��*�3L����ֲ��G�M��;۽Q5z8�a��q`]����2�WFt#~��+qjǞ����A��n
4�*����E���@�%��"�«����ز��� 3��I��߉P&�F�5zm����"��^������D&~��u������c�9J_�H��4��E��>l�ԢP�o!FMaK�+H�U�S�����A�.X�{R
��(��N�zl�#-ۓ���^�K�?�T��Pě��t������H��޺�e�i����lOt����.�7t��������Ơ�~��<?1cC^RQ	>��_�-�x�b�n��M�K���L�%m��Uç����J�k�!/q����7��gnW�
���)�����>[��2����i�x�P�-��H4_�G�^
;�f��e9e:� p݆A�v�ӯ������K����qN|�V|��z���y���0%R ������-�/'D�R��JZ�+�0��F#�Y�c~Xk�f�K��E�.9��_"�ͬU���c���\�`q�	��F�}���^t���ӏ�z�J۲���4+S _#�@NaEn¡ma��0R�7�Ő��[���9�CZ'P��cد/��`aX�I�h.������Ԃ�ɻ�����\ICvѹ?�#6���V-^Քt���a~�M�y���V����V�H��:zo���Y�+z��9i?+�'O�媢6#oT~���CObu���>�
���q��6P�HF�����p���J�X9�Yo�N��L]���H�D��w~&���	H�����R�oC����n���9L��7���&�j+"������e�ȥ
�E\xYа 3J(u���t"��0��.Ka)�rr�(�l��dj�"��������%#�����l{T�ˉQ�m���ax�JK��1��������Ӊ�1.C��8�	y~���9�ԢU�	��}I^`A�dD�㽵�,+w�45e�Y�~z}����S��KbTJ���r��ΏMI���@/��X�U�-=�����^��u���͆�����&I@j�A��np�gԸ�˛�]��Uћ�}\#�f����sa�)���R[���A�N����!�C`���`�i���E FB�˝�+��Xk�c���w�QW�y�꣢)��hnn��<����S�JO�e���Ɵ�&!��iT�nġ��_N�R�lY��@P$/H\8�¸�P68�~H��,�jڋ�;����?��E�R�y6�䟈��yP� 0��1�Q�?T�~��� �Q<`���ʊӻ��D�|��~�1e�z�o"��W|�%�/Ï��N�.*�b�m�Č�)�.��u�	d��%��z�<~Ul�#� *�4�l�d��.�w*t�z_�np���.�U?DN�u�7��IS�V�9��֐e���Y^�������������T�hRԺ���3�/|�%�v ����*��7| ��r:���rV-�f���DB�����}�
�	4-�|@#��"Zq����j���ɥ���p��D���۩�^{���ｼ��쫗�c7"�?�<�/A&���G >22�#�9e�)���b��&�;�~#7wА�d��_T1��(�)����y�z	y����W�rN�\�~>���8��H��0���g"�g���,�NWi7 �u;t�2 �ƍ6�ac	��// k��^qb�sG=�՛�`�����va@�I�-�3�fw�U�ݽ1�[/_��3g��d�M�� �k���)[������^!��\��G@���n��jʴ�w�N����,Z�U��]t0�<����f���/���T��?�n=Sf�h�.�=�m�6�d�yoa�����X�?�('����{��kT�)/�|�1�P�5�S�Mz��-��ǵ�7$�b}x妞�������y�.T�6�3���v��,ټ ���
��$p901|�gs�8��_���(���<�y��LlI�����ljj7��橈�:�x,Y�<�Ƌ�1U�2=Y�q�3�����%S��OJݳ�ug�B�ę�2�4��K8%�GЪ*	��У	`����b�֥a�0�h�a7ac�Ku�5
����)4��5èN}��I���;]"2����iT�Φ����z�I���]���0�w��i
�ЕGS�&���4�����ߟ�l��i�i�XC��i�S&1ś��h6��S 5�Kѱ��[�N���տCgQ��2דC 8ª	
����!&�+�7��V[��\T�ۥ��/�i`���<��俎��T(Ga�5�!7�����e
����7ä"K�1���GLPԝ�n���K�	T
rV
�E�xzZ���y�����r{M��T��<�|9{�}<UY+�T�����lz�Y`Qc^x���R��<ۣ ���*��a.!� ��FH���$)uh�/?���Ǐ�>ET���-�-I8z��w��}���-���pJ�l�/5�-Cb����W,�#�;��GS���X	����.�px,">h�_g1t�+i�Z��,���� �!P*%��	g�=�t'#�X��Q�����e[�U���O����B�����Ur����>ǝٶ�,K�.�h�,�b	>���|��7"�ۃ��k*���xw����<gS�}u5C)ёwl�`b�6�~���Kn7��Y�~c3�Wmxd}_l\��-��2�m���h=��E��u��t�^&|��{�?��)=	���S��Q��y0�c��"��F�#~KT;?fӟd���*�$�j��q����ަ�j҂T]/ x�n���x�V(p�F�"��c�x�J�E4d��M���Sőz�MB�*�"� x�oeE��%�%��n�T�t@�̒�߽H�c���	�=���\G�2R�ߙ�N݉(��t��u@2YD��hXI �N�S/ު�v���� -�_�˕8S�4i��}I��N����_t��l��?�����Hd�U��	N��7{Ƨ��=fx�f�C�͎�;nF��6n�M޼�o�J\_��h��}�އ�6BQ��׌�jx����ː��c�w�f �xU���H(����&�E����`�k��������X�˯}�@�.Z>]��@ؽe�� W���d����R�'S@4��c��T�}�0M�ո,�wEC��YG�۸�7l��{�i�pyġ�Ba7=��p�1m]	ݟT��>���QvD��J����l~�ρ�]��,z���*!�q��əIq���w�q�h�h�i����+�+��w���A����E5���n�5�*Q��x����� ��A��'N�YNs&�}=���8�����m�/s,���a-G�CZPW L6���`�0X��eԅg�B�\�o^@�t�蟴��MU��/ǝz`u�O�U˂��������N0���%\\L{���Ձ����� ݴ�dA��U����QZ	�{�"ImhЌ��ٮ}�O�GB�s����?��^~Ő���/��@��A���d�{�fҮ��(�nn5�6�.�����1�J5k�����P�[L�ZS#����ѐʯCs�