��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%�ח�.4[s���4)�9ђX�~0u�B�(���|+sP8�D�mp����
�=Dv�T�);z�G�z�O��9-+�uW�A�0�5��ֺ�H����o����Xq�SA�J�F�B�e���"�:[�1����1uj�	C /�ŀ�S�U�2O�:����UH�@>���-��:��Tk��0�������YS�q9{�S�Z�&�:z�`�Y�� �n��J��h_�8�G�pU�s���p*���H�Jy/Wu	��k�&���:_��M�c��N�ZZ�K�����U܀ZE:�?�m�q��ʒW�x�1����P}��-S̿@�ts7	E���$7���&�c���9�:�ڋ��Y}�1�����5L��-��s�pI�&�B7bq��&�� B�R[Ɲ�C�:�t��<F�:�����x��K
�O���"ճ��5-��^-I�I�G�T���.��̉5��$���2�O�7W��
S������^��)�5{d�RdՈך���$=�<|�;�E��)����^1(�Wq@���r�)���Γ�NW�+X);{�S�� ��������:���x�4�z&�&R��KQ
�S��y0��-)0��YX_�=�Q�]Cf�[��IP�UUX�7����D͋q���d5�m��N�I]�S���M���ز^}r������w���)K?�x1�]�P�I�Y�ߜ��y�$JX�2�#��JxD��Ս���4�=�L�k��ǘ
!�T��i�)� O�f�yV0t��'�u��=#*�{��2~~X�|��/OL��j��"�//ċ|��2]��c�y;0ʋd�+贛jr��4��i\~{��@���"�K]"�����2E$T9!Fʐ��U+������{n�tJ`��e퉟�[s��,����}2$���,n��e��#/�Kʧ�J"7��Z��`EB�^�tj2��9�ٖ��K�(4��g碥N`���/�>�⹣���i�*���H$�IwU<�웇Y��h�!��Z#���1b��a�����+#�NB���H�����Cj���vq
/�0�P &�l[a~5<E@��~7r(3/��.
9�_mM��z����G�4q�F���0�G�T)GҠt���Q]}ݠ�b��5ʖ�޵N�\�j��Q���G��w4�!Q�`��+�t9;/��Z6AR� �?���Mm�J�sJRڕ���lۖYPΈ�Yw�����'	�LԵ6����"�Y����u=��xE���>9|�B,���!�?�v?R���]i �O�;�������=�?������7$�t֑3�S��%���Q\l����-wO�5�Mk��:����t��l!��.��N�����~��O��_ ��l���n�i���p��ʎ��+�J`�����t�r��+݃׈��j7�n���a�Mq��ק`��Z����)�8~��T+���������[q6m����M�At���k�@k�E�_FST	8��n�V(�l�4y�"IKq%+z��0�����F�������J��t��$-��Y�i��['qW/(��V�@d/�8Cga,u��x�lA���Ftr75�XT�L�ͭ�%ɂ��D��+s�L�R���ѿNX6�q���4�����n^֩rN�t�X��أ�햴B���1�
I� {��!��@���'�% ��.��Tx$��E�P�}H�������c2'}~���z�Z��]TbS`M��eu����r�W��ip" z�|Zd}z1=J��.q��%�e�l�A1yV6+��
�ى���9P��|��H�w{�����"����.�(��1���c�m�5>�b��Ut@+����ۣ�?ɩ=
4�
�l{#!-.i��5c�
GY�RR<fN��ސі�Hk���瀯���{Z��� 1�`�L4?F���c��<�{���c��$�5�Jn�ȴ�N��Mf��:O���eڗ�w��>�$�@cMoJ%���]tT�aݲ�`�U�r�~�=�9?����\�40�n��K�²��}����/��?)�=��ߠ�`�1�\��#�璾��C�F)���M�:v ga�0��>폿����D|3�cR�T�@A"Py#�:�%aէ@�O<O�����re	i�N���sܐ��5X6�*8f�W�h���oB>������P�����jV���Pي��w8����c!J�x��P��,��]C��hM�8�}ޚʯO���t�HK��(f��U�n|�����'M_%/yXC�p�����C�ߌ̷h��k��#�.����:C�3JUN@}I �H��,f�
 �Gi���j�$�o�鉖}(�虁�����)	��I��/�Z]�t����Q�	��p� �|-�<.0}�y�"�ǃ�� 9=���~Ҍ�9buQ�������a����&!��"�L�����
o�ԓ#�I%���N�$���tqZ2�>�A�6��~,���9!X¥�/b�nS���	���BF�Q�i�f��:>\g�!��0{��P��-��k��@���P	�����o@�� �rv�h�h�*��`�����>����EW�6L�t�4�H\s:G믌��ؕR����%�:��$�,��dgY %����[.'7M�̘�Eq���Nc�<�ݻS�Sԛ���6X�3�*��j�:�A���۲`�b�3��t�{��tC��COVj怠Ƭt�-�U���WDv��H�v�g������(��*�E���C�>��q��7����w�m+v1��TL�t��u�)4_�Q�j_]I:�C ���+��)g�0{�8s�{��_��W���GӲ�{rd|;oU��G�p�?%{g�6~)n�#��� ����|"}H��[$1s��-�&4B�aƮ{e������u��sJ�xؗe��	�dZ��BY �V���Չ��En�o��k?A4�!6�C�$FW�3�r���eIa��I���ߣ�����l]+�]9������I&�:r�?�/`JFe�� b�J�SFy.-Kv8T�-*��� -5K6b��6˯رp��з.<�=�_N4�&󛘾�CYD�F�k��a���~�����0�����&�k0PfJ�B\�o�p�͎P[��=
�rXw&�}��^�֒ZR+�J�h��8�kW�h�Ro���^M��UA�X�<w�V?��)ؖ2b��9�	������X�	�N��f+�1�@l�
P��Ê�B���r�Ł���~T�ឱk�5���M�I�Ffxu{Ly�t���ӬN��0��qIzxX-����*���2��8�#u:��ơ^]Cd	p�����(*s�F�).B#��� h1çMh�Xy[��H�U.��Z�G��5�R�!��X���
g#y�=i��n��hQ�#̝��v������86��S:�C����5�P�����-6WxP�5�v�x/|(��W��膈���&G�����A�]���o���B�p�I����h��;�m��V�q���^�9�i��ى� �]txqHT�D-�Q��9�}�dZ��J�y� ��#'� ��-�7�)���z� �����]��ς�C;f���_����!:�V�� �1�>:�ŷ.�v���\>
'�1wOá5��gfb�'ő��� �-Bw^5;�3�L�Uu�O�a_��sqr�Ɂ��$?��I��WjA�����N��`���RA��.V}.��W�+�ЋH8]��GD��t1�#ćG��$תG����R���� ��ߑD��c�>��E��E.�W���'�-��p���M�]�9`��4 c?9z�˵ȩ�Z�"��T�G�X��	�� =���_�_�!^�Q��Q�s�KH�/eo1?'��ڷ��,.�T<ܯ^�<��$x����хJ�Lu4A&F�i��Q31Ň�I�}�b���.{ϡ�8�s�]���_;Ř�>��'��DcZǖ�c�!��xD�]́"����X���|F+�w���
�4�Q������G���6��-�ą�[���1d�6��ߥ=�5,�a�+� ndT_)�	�O�"`���UP�-3_{�9{Zy� x������VKz�B�6��t�Y�x��ruDH�S�ʶ�����M��ߚ�d��h���i[�ptB>�{�P@uB��v�HNߔ���E���#��.1͜T`$!�� .�͸ v�����������R8��"���X�%��I�8gZ�#d�Tn�"⧴�\��;Io��9���:��H���ǁ��IJԎ�#f]��K*ߛ,��,kє��9H8����I7��Fl�({_�$�8F�E3T��ym9���CP�lr�$s���+6�)����96M-k�2�'�{A4��=1ӎ����Z%�~W�sķ���*X�UC ��� K��U��'��:�b�6?�澹⊚������v�#="�G�t�h8_%�Zk���3E�݁���l��$�v�����
U8L�k ,�R�����k�?��(�;H�����ֹ?'%�[��6�������]��=�(�t��i�sŭD�~�'f�[`���ÖT]ȣ�ܠr��7�	u1�ζ�����M���2(����XO�)�Vj��JE_��������^��|<*�4	\�-S� (XيU��#l3��x������Q�:�=7�
yv�Ȕ7=�Vs��I���Ĺl���4�_��@nsp�G�e�O������=d�_��������yv�gZL��|���)Qxp��.�����M$v�w�,+I�.�K�|���C��?+�����=�j���M���-�׆��Za�Ѕ�^������j����q��8���39B�7��&����?�X��).��b�*_��.U��1�?s�rN3&c�_�>n4)��}w�#���2k��L�Y��F�8���ii�`����[��ey�2@>�4mr�UrD�3'�u�H�n�;;V��Og���0v�`Q�9���5��t�'=���[T���߷b��~Q��a8��.<��rJYb�O��#0��PsZ��E�&��N����8�Åk��p��aG�R.r�W��NOE�h�~]��=��y�0~N��xY����|�J���0���꺡�+X��|Ǣw.tH��#^Ԍ�O�<���K�*�ymC^(���8d�nk̓#�<#�Zy��q���M 9��\0nkn���৓���#�[�JV?�tJ��h)�Ɉ�{��D��>eI��q�qB����HbI;�,*Ǡ����*�ֈ*�ݪ���+�_k�p��5f(5P��\x�Y� ��[��&2�!�=hm��<��uf'��������E�ʇ@d���V��8K����lTW�y�2A��'u����'��J`�;`�؎Ga��K_/��SD+f2�"U�8n'�x��'�g:R]<��ۏz�H���ϵ)6e���E�F�I���ME�֟Y�-��4���g�Up޿�J��;\�3��J��"&����>u��*9����f�- �<�|�P{���ft�iy���#Ϸ3���
��K�f O�W�=��� ��l�&ځ���|E]H����t��I�80k�58��)ms~��p�.��@������m;Ȝ�E+L�ʅgl�O���U��6��ȧ ��i���7ơ��)I�k;��@�ԫ_�MH]�ϻx�����ňH���~<�К�uf�D<p2X#b3����̙���yBo��l驍>���ХV�<u�v��)��D=oΤM�l;��+��ϛ�JT���S Sd��)�f�o��(>�WH�*������-K� ��c_�����*���y��VM�狽;��0Y�³�sG������'��Q��â��9������(n��Y�������Ϙ|��D�d�mr���$8d"N��x�j�"pO��?�4�=g���A�E��tAU�xF�g�sw���k]b�%P���O���&Y�9j��gBz�$�JST�=��|0P�⥍+��&�o�1?�P$%��F�@���+�/�M �+W�R��Nw�����/8yS zo��;��u.���0Z|�ncm�-�����헜�{S]&��X��J�H�L���p DvzR;�?�Z�
=E��T��I�sQe�)޹�_2��<d�`u�3��z1���L��d8��	��|���\e9_BhW�ɯ��TZh�[f_��ݽ|;�Lﶧ��9ā��%���-���h��1�%�x�`�5�u��ОX9��J���(�,ȁ����`��	�3h�"g���q_��o<��`��#�w�8�3�C�h�ȝ�巺R�0.��B���ە鋮M]׋Gx���>��t*��౎�V]���]Ύ��uX�̛p�}s�.�,��V��Y4�L�!��	x���[�n�xuFs��O���IϢ�ʺG�k���Bg~�l�3��k�ɂ ��mDV's(��A� S.�wG���ݔ��O'Ȃ�$�m�(b����xz��q��*����;�JN�vҹ�,Җt����o�j��4e@p�/2x<\��b/A��`��3v�@)�_�:o�B���J��>'4�>+�Y��t���;p�y4u��(ƅ�ؠ:=WV P�����$x(T�K�.p�@nb^-r��q���B��u�������Fm��m�oN�ƃ����+	�����9G��YEը�f/+8`m¿wN�p�?8�2���v|,ƪ���\?j�n�of�G���~\Uϖh�@��S��in�V��Ȝ¸�`�/OGo�Fíaf��NF�������V���2Ó�(�hJ����s�ߐ\�r�V��F
sAv5b˯�&���,=��t�*�z:��ܟ1ǜwtF��a��wHlR2)�V�u���柒Ag�!1�� H_i'�URÚ�bَ�;�����M�R�8Vե_���ۃu��?j-h�N޲����/?RY��b�Ml}^��װ���Ҵ�(�>��%�/����I�T��*�L�L,�H�.�=�p�l�D���!0^�Q��Ǵ%EX��\� �gT�:�0�bt	�o�n���7;!m�q�����<��5���5��'n�x��ڭs@3��l�x���B:��O�a6<}��x��P@���-�Ys��2��H~$�GH����@\��$H5�:Z�H�E�}��r�� @�8��1�m�2 F��F|@]�)NI��q*3����Z��E@N��$@th�	�=�i['�j�G��1Ahl��`�ښ�8P��HꪆC���C�b��a��a,L�����k���MP�jY��Y3��OM����+���{��?�!z��"+b�����v)�������{S4���Yc6���F1���-&�3���T��y�>�w�EB�I]��@���m�g�ZOV4�VW)��JRA��%�Uv;C��i��(��r��l�+ m:��a*`�qY=R̔
�~��`��3ҫ��?f�>��=�+�Ҷᐠl�3���-a��Ъ��r#�O���S�p8A��T�5�>�m�^�
i�oh��G���*��L�Bj95�l[-��FAo	��`U�����=(��8�����%�[f���ڦc��ᣊ�@�tXB]��Tp��%��������[�Q�~7怇L�+�ֿQ_�_
N��j��Ǻ�rpB���F�y9�j$R���\A�Z�����۫��S���G����	3�n�}�쬁*�/�(qd<σbF%W��^yy��J�E9���I�:��U����'i�U;n��\�D�P�:���������%u�m����H��>���,_D���)+����iV1OΎ�h��`�[����pp7�Pj��+w�\g��H 9Q
, �lQ!�}��_���S�\���N2��K�V\�!q���Q����lK��5I-٘Զ��%Jk�r5%���-�"j�1R�},a��o�n�ہ��Zo�ڜ�^�v�J��DR�֩�����Z�Wbf��q�z���N��{Ҥ���$�m�ĸ<����:�/�=��4����G��$Z����A��Ȋ�T����m��(X a�ҥ/�X����g���:(�qx���JL̕%��ݿOL�mo�T}��ƴԩ�vLI��M�6*��M�сM���\b��f8h�g�n4r�ON�?�`�N�q�?�����i�"T� ��%�^rۼq�a����a��������g�&Nx�?����������j���=FN1��o/�����z�(=�7�|�����#j�=��;�Q{���Cn*���u���hQ'3�B��Y�V�k�xvge���|���5�ܳ�EY(��]5GRۤ����I:R�FǓ�|�-��f��R�QwY<�S�y�d�.랖�m�� �:�M`�T�Q��{F^�����-JiE�dQ�E�W�i�z�C�hE��~�������rS���>��r�����q���\�jI�i=�Ӝ+��J��n�_�[ȫKγ؃NU���vU�tحK�����Tb�	fR^��7_�c>�R�M)�M���E�8���)�h�����tP:1�K�y���V��8���a��q����Aڙg%C���G�3����Y�d:-�0�s��XC�w71/���1!�W��'{[Yq�XL4� ���Y	Y9��<�gY/2���̦֥	*�e�V,��N?nc��]��B�wTh(/�/;�F�>�����ƝJ+��G�62	s й7�����R�?"R-9�a���dΛ�,\�i���6�\���D����+\�TinGf%mH}S���f�;n�����z_ܴt�r����|������r�-�^Y�棉D$��H}�㯠�[�W�=�0�/�񫣡 F�J:��1#*['�|k�ok��P�	C��F���Q0�8B�C�d��}����sLY5D� '�S��K�Q��®dm
G��~��T�W4{h[Uī��G��t�P3C,5mM������W`\��{�pS�����d����;T%��E�+w� �k]�/֚��Ҁ��_��!V-F��&��-�e*-�^K�ryRo4id���;��q��:��9|�����t���5�S�Z������!�΋�t���*�ͅDMU�� y2��g{��"{���5[kN�n�0����Q�B�d3��^x�#�����p9u�ѭѧ*�5�+���#5�l1�5ߐ(`����Z���֭�A�I�w��d&� �B�3eYY�4-���������K���3 �	�@���^�62�%�5R����6ǕX #t�,���x��ګ���z1�Kg������=$����	SQ)|����J7�4�;���3� ���~���q�פ\�kK�������-t%=�EՐ[�'W�%�	�3k�7Dy2\��Jr�)����U�(9�9��-���t�+�&9T�Tco��<	��q�Z6N�}a�$-u+wJ�s;�V���EB�zs/ԗFH�������d�����`��gt,�A3'z�YE��W�'kπ������8Jd�	���.q�Q>�x����bpN�[����6z��/�9������zn�mځ�������=o��>>����b�����^ށ��t�|��+Y�����k�\3��'���Y�F6�E�>@��Bo~se��%uԐ�J�_��o^�*L����%m/����h'�'���
��Ѥ4F:A�Mb��~E(I�w���:���$7�T~ݙ�k2�R#�Ք����w|r�yV�'���!pT���;J)!�����C�P�]˧hH�M��k�o�
�z�{l,{��A o׽��������=^�om�E����IO6d�rE-����SDD="�W9-�H�Vm~�����'x��=&�GC�B�(\�/�)e����2�>�F'ʲOȢH��3�T�@�:Tb�w�fU�bu�v������y:�KUj�O-OG7���[��HY^�	/�j��u3Ҧdoe�o���>5�3�"&�}��/���rA�oN<�ӑV@$�ă�݄ Ѿ�H�y����X��p���Cޟ����S+���BM�*J鄜ś�,j�D��`k��3�'7`��	�䨔�.h>�_��B�%�*b�Q�ݿ�8 ��q+��Î�W��T|B��������a$4�:^���'�6�xf�@�P��҄�ģ'��d�N6k��s��.Vr փ��1�<�*/�J���<:_�4�{eJz�767f2Z�]˗Ũ���)A�h��
���h'�U���.���1Nyq���陖v�4������w���ơ��<���@d&�A�'��$��4�A ���B�vVg����W��
*]���ط��+: 5�Xݷ���A����x���mH��BL�h��M3��)�*���)r'7���A����dz�����)�j���_#@�pk���2���Е�T���H�⾍�C8�Q�_����"����5>�A��؏��]T\�z;!AԢV�{�L.ل�8㿚ι��F�-�3(^�í��B�\�aN��Rmg� ���L���G�&�vu
��I�-��J.�E��l2 ���ɴ?�w$[M4%Ӿ�Z�"�#~���B\�iQ�s�3V�Q�x�E[#L�?���g`�pg��[�ћ�D���<Ӟ���9���c��kE�4��-�_���>��ʍ�хb�ڎH�+Сd��d�:c3�v�s" k��([S��SO�M�\����qM(����u�2Xf5]_PU
et�_[۬M�pb`�T�١ilZy=�,�������
�jW�3�"M|�rX�?68�7M�#0����S��x�������y\���h��wJ�~๤C�ԩ�iN��Uj���`g��S$Z��ƭ���.��ޙJ� l������������2�S��rk�/Jw�[TZ:7��3�� rd݀i졓����O�l��}��O�I�0+�� �c�	�U��#�"J���A�C���͎㚹�;�z�$��a�6$���a�q� ���xtQ���K>U8��� �B�Fi��k2-{|Y���Xʼ�w�oe�|�>� �V ��@� >e[�_��q�_Qr���+u�S����-G*ϱ	�'�d�\�i%"�a�)
ͱ���=іi�j[Ȭ�B��s�
�_��$���_��JZ*=�0�yE�#�>�n+�[̟�W����8EtH�U��N�A���d�c'QYJ"-��v[tF�䗘���#��۷��a�>���#�W�'G�<�����.z�J8gS�f��?���A:�t�ˌ�G���nS�& C��گx�	���k���L�|��O$��U�#`�T-Oe腏V������>�Xk �7�#Y��|��E#�gp�\?����Cs�ǰ�s�e��FY%�����_Y�4���W�O�:oc�>)�>$ΛH�px���;Y�|�-���Ǔݣ��X �@^ݝq�c����;&��3�lk�D�����_T�9*.N�dbH��"�Z��=��hP���q�G)$�o�Q�cl�b�r7K���˨�8�3����x�7)Ev��Q�|���:Q�8�us��=�E֢�ccb6t�bB�Lє����ج�W%�h�A��"��|��C,v�벗�z>S���x�.wHu@�.�
���b<wV��n��.x/,f3i���laa��@Ҩ��1��Q'�ο�q�5���;�:�Ӕ��pM�c8���@�H�#@[�A`=Ea�a��p`:R�3� Y�p�&�2mE����TG4̝���������,6���Yݽ�)	2�H'q�i���*NP-�ppYg��D���M���T�rqb�6oX���[�&M��%h���qb�O���8�CF�p%������d�o�~=ee���w�"d��T %�+\��#���}�xK��(��Ya��4�:�b �����]����9�.`n�el�#��a��{9���2�`����t�+U�Y~q���ػ��ё��%i-E6�S�ڷ"�=�F���t�jă<�Ih�.bc.��p�[�'V�<G�ߠ61������ss�Z1����0���cl����K״hA7�c��e�8�nOxi�cl�fXmv����� �B	��-޿L�*��}�r�a�^�sP_�CO�,�$� �X_��� �S�8T�/�_��ݜ�w�����KX�������h�hĞ��*�ZP��7qu�.7@�L�6��"����K��YE"~"�-7�:E��kX�4���S8` ��NU�*!����6�?-3ԟ��1,l��ޣw�kVΩ2\�&�X�C�-��mx�Ow��J�0�4��d�O���{`nIg����y>��؎�$ɍiږ����a�5�CV4�F�G҂?�p�푾2�����:A%e;����׋��g��E+<tA}_ņ��p�[P��p
<���RHK�=���n[3��{�x�e5�~�qv�	��}�8\������;q刱t�Ҫ2���0^�d"���xڪ"kLΝ,0��c�D��̝!fl��)�\!��4kw�t�*W�h��*�V޸.����E��\�)B��md������mm��M�����%��_����E���z\Ĕ��_vX��,�K��f�f# zz�m"]�F�51<��sM��3\���/R����Z�ʺNZ2�Wb�H9C�(7����t��g-���|����ֲ"���+T=MS���3 �7�� ��2?�*˙��~e�G�
��j�y�1��ƣ#��Rum��,@����o���V_jA4�?��[0�u.�0�iYrN�����)�3�;>�wr)թ���*�OF@\���a��,�R��0w��g�)�1d|�O���3}�{L	��
bġ:��v@'��>�if�ug�p��C�İ"��꺎DaK����mM61��ov�<���=��QOla�#�`�	s&��D�������1�,��ڰ{��y�j���/��J�4<�`���[����,�U��Taj�QuV"�_�N$t�:��㠗/��3/�zًQ�;=<�O�-���	�j�U����1.�ks��T��鯁���WG�e	�0��Ɍ��1�*�G������C���jn�i7�N������Sӂ%i�Ы�Q	#��8`	̝�a�^օ\%��,�
i%h�g㔓P,��qЖ��^��F�?�u���T0��@�[0t�3�>0�\5��%����4Z9�a1�k�Wp��ˑƅ	�u���2�,Wr�A�[�Y,�p;��9�}����x}X���	SX����ߌ��<~aq���\��w8��6f������ZmB�3�1�f�p����E~)�r��x0������_ �tƔ���	\��/bET��ꀺh�������OLպoY��U��<�$�m)QwB#����&�]4Q$��imԑ��m���|���m�Cd��]��SS��fP/ua?z�����S�/Z���JV�y��{(�]�FK�~�"�`<��;ǔ�dXƆ�k�cSh�w��[i�WĜ�Y�A�լ�G;�vv.�)���k �zp�ɶ'dI �L`��7����A���f�(�:�Z�� @���q:�0��K��9���"��̓��v�a�c�`^�yy`��RN�Š`��7��ߟ��3uԱ��Y^h-�U���9��i
�$�Bf ����m<e;'�VhHc�͐�<�R?�s�,b,X�
�Z��N�4�&-b��Ӓ��[r�<I��q������=��[��j����HF�Q�rv��j��C�� � ���j��N�Ԕn7mv���|?K�ZD���'�-}-�l���*���ʃ~�Lx�Eu��
�I�W�u�PV+_���ɟI�����h�uiI|Y�U��Ab����߆'i����sIRuZ�8����ջ�Z���:_3o�����i�_�'��� &������o�(p�C�����b`���n~&�kC?Iäw��kRf5�җ�������%�\ﵡ�E��.ѵ��4[#��+F���%�dY)�HS{�����2��47 :qО�%e3}�i"��o���~N��D����8����NMB�g^{���p`%XҎ2J��߽-6i�{���6���;�C��G���Ie��[�ӭ��)P��M$"
C�������bV�"*���"X�}_�O�f;��́;���٨ǸĀk��D@�>��vlq�7��{@�@�ԬO��A:� n��������r��L(j�A�zE"�pMڽ�D~���x��8���6�i�~4|�i���b��E&�t��.a�"�I�ٯ�4P��B��Ԁ�!���X����`��������Ipx�E(�~hӍ{���C�@u16d�aw����M��_���D��9uvD��'Q&0#y���2;E[�Z�/��>�m���-�����q����l�����k=A�HXNU���72���)T��
�i �Q���w�3Y���˗n�Z�ے���gO�������L�0T�Y��l1���8�ф�C:L��QlbB�<�-�A�>aJ7�7{QF���%�"��,��w�./�,M�"�M���2��p����UN��o����sKǜ9�iq/P
���	��X(FK]�����2�������ّ�O���˗f��b�B��	c�q�d��Ss:M�잻�J)�O�rQ�:o�8���ϵ1-�8�~�z'8 m�����5����x�b])�^_�~@S�a���8��0�K����h�y�[<F�"�l@n��E��m�)�3LU��Zr˲�@"����I�<Ȃ+a�&�u�\��?܃C�)����LQ&`����*x|���v��gU��Eе�r�Mj� (&p�1�ʭ�d��َ��� ���I_�~3t������6�uYIЂ��J�f��\1yt�z}����XV�(4��wcכ��:1�)G�J��v��W�wN:^��[+kx9�Yz$�e��5�x�UN`�B��.zo��e���R���5�f�f5e��TA�"~���ߴ�������}m���xb{�l���0��#�L�|f����HԆaJ
P�~x�­%g� ��`�9�C&���Z�[4�k��h���ڧ� ��K��B9�k�C�����^-�~���QL�ӡ���N.��"M/tzڱ��d'��	��QsQI�!&R�����l��{�^��Әq�Q�PL��!i���H��V� ��L񡟱m�5)�(:.�s�-X[��mڶ��E�Zu�ę��:
��sTM�7e�@��E�w�n(�9����k�,�l�UA�@ۛI��UV��$BW"�ަ���~��	��r��lD��r'r���|%^Zxm	o��@�̡+������˴OU-2��d�^�u��H�� l�^wI��l��DZ�W�-9�)K�lJT��]�0�N�`�B�Z� x�s��h9�&��4�h����ܟDJ+��Ⱦ��PX����?�F0�8���$�9����ēE�}v=Pu�y|0���~�Kj=���w�^p��$b��QΩ�9����E�=r�؏u۞�B��Z�0eO^���E�&�0�$�M��=�2LK���.z��2�;��6���f�Ml��7�G����ja�mXf4�{9�(�[��Pĸ[�������O`N�{w�4[�ר#m�[2�����v���Z�
��&���1J��a%�x�	����pE�&"����Kp,�{"���x�EK��Z(ZZi6r�[k��F,�D�1�����RUsȵ��e�e_�(�&>��!���&�a�͒7�l���B����;�C�"�^�RLV@����_E#yag���p�J����s	��ϢJW��]{E'�Q��b8�k�Owh�b2uC��im)��D|���;�D��aX�d��X�%R��M�|����?����!�4�vo���5"c)�UH����AN����}�>���V��&�`o>�����%�dɄ���Õ��wET� �øV���DX�UE�pdyT��9�������=�FHI����3�|�n�bd��Y���KP���]%#Ѻ�[v�ؑ+m9�P��0�.����Z��^�?��:E:eh{��v�w�����K=�M�2��R��F��3��D!.Ƣ��YM��?��o�e�EMf�18r��n���@�Y�O���>��X���3)�7uN�#`Bq�Kn���bv��9������<!8��5��7\4�C�����x�r7����t���|��c�����n=�-�AH���>l�«Pe��2"�
��8.|�s߄��G0� �;Ia��kS~DUy��pِ�f&�p�eU�{��3���5��1�EH����m�D��8��K��SIb<.�'�q�#�U�{��B����ka���HRb\��|N����{l��d��cA����JT{�<{lш��}n_ �$��k(#2C&�&������1���c�T7f�4FA@�aC�$G�_�e ˎ%�Cz�i-�Ŋ;�o��?��^�U{bXM=�j7����U��Q�
��,���/u�B�Y�ei�b�U����:�0��D��H#R�R�)����҄�����=C��*�W�/�k>�H틲�����[��#<�a:���y;�ɸ��b`������7�����m-�������W%�H�~^�s��	�;Z*|W�M�Y�F�����wϧY_�Z+V�V�}yZ�X��$7&���2�$��~kQyٴ�KBs\�B��6���{�"����y�:o�gq�qP�oV�Y�Y�q�˥}�@��IB�Tb�1�fu�u���~؍m�wyA��fBѷ(*9.�}V_R�t��dj���M	N��,6��)0t�~�Vȇ�B� ��٩��/���F��g�x
6QLf����x�C��Ɍ��z�h$�Q��fA!��[W�����M��h�ƒ-��?&�F[�j�~'�0l�o6�P/����hU�J�rh��.�C��,��&ޛ�ć)E�;�(��������,�i��\�(���Q�$_O �cuG�B<��M��q7U��b�v�\���ʆ��#��m���s�B�E�k4*h���ɕ�0��_7���gV\�Q�mђ/j N)%�!Ԍ��aL��U��t�D�;��K�2�ݎv\xIŔ��ȭ#o
���6 �$�b�� 2 ��=�Z�j o�}O�TJH�ljgF)2m���	��e�3^hK�����l�C��[�x@������>�%%[תXNk��+=�5ڒ ^�H�Ǡ[�_;9�R���P��o����� M�ȗ����e��:�-�J�9�i�gOP�P�Խ�g�-�s�ʓ��d�ΟsQꜶ^���!B�t�{��M��,QQ�A�a���������J�l�.�]ç�9|i�V{�]Qb�z�r�hl{q�:�f�����XK"��0t8n�3�(u+^v��&/٧�a�WG<����H� `~������f���;E��%��b\BHp!B�L0_�� ����o�Q�ģx|!T�67|_�p��ݣ�r�厗u��I+��W�`��N��*��m�R��12!�B 	Z�����"_�<yf[-{�&x$_0U��=���j͡���l��2�2;��[��6f�̤��g!Pa�cÐl��>\ v6��{2�4�k$P^�H�c-��-b��xZSgw
���<M�>^6h-���#k�k�� ��
O����u�yٖ�ٻ��ej�M�
zP���tS-/ӈђI�<;��B�lʛv�?��k̞8Ai$b��#��^�B�W�6�c��� ��h�78��v�`"�|(q����rs .��#f�́$��(!n���v2�޵e\J��y�)�5¹�����p�=﫪Վ�[]���n�nD�t�N�ջF�0,[�����bFF���q!���$ ����c�P[��hO�Af�Ъ���SER�+5�ѯ]�A�"�G�vQ�)<�B���V�9�����`��Eʛ�M{�-ɂ�� ���W4��O�h�X4�Id��b9;��tn3㰾܆P8�j����ů��p�	��>�4*����?�GB�и$y��q����i�a�^�؈@������5_5A�X��,��s"�@K<�_y���G�h2mK�^[�Y%l�nP�V�
�B1�aձ��VZR�p�4���Yd�����Z���V����]�����F�6C��.�d?����0��q<�F��2C�40OGG�f@�AG�SZO2Y�h`���2Ô(i��������/Px�r�AQ*�t:P�o�z��6JN ��O ��� j���{��NB���A��	c��wXiE��Z�.�G�ʦĳ\k�It�j���W�F�� 	�3zg!��:�)N�X�Ľ2^u0"�����K�L�m�=�և���V뮊��]�Sh��h��U㐮P{A>�k͔��Y`* �y�%����3��&-���2�Pc��z�b��@�c�%$��):����\�D2˽.*Xs��w���u���-[(�1��X�����{C��3,�w�}F;=��~%ۖ��2��	n�f���c(C7�Ϧ�`��15� bxI}Q����yP �)�5⥺�
�]�	_�g�@�9�Vʭ7��O���/!LC��5(���1g"l%2�Bӑ
.�,�oe�#t^$��	�+�-�i|Mᓄ��F�n�Bgp�^B���B���#��=x�܈_�����E�!
��N�w���C^� ��h�����ɔ�\R#b���;�c��B�E�0wM�!�`DC7�s����}s��8,�M[K����K`�����S9�6�Y�,��2�|��0��J�(����Z�e�c��W��L��W���ck��r���%x��q������Xs�ĤQp��-�k�K�
g���o!�qhQ_BN��>~��[M�7��e+�JQVXHNn���,>��J���Y ꆜ�2�εo��V�jVTB�T;���-Ѧ��(I~҅C�©y���P���&������-5'�r������1�I�l�7�"���H��mQ@)c�!vA��;�[�j�֐H�`����������L�\~P�`5:���d���1���}�j���I�!�Ihb~`}▎�Z��/������ �ۮ���Ȕ=��;�]HG�1�c�,T�j�ٰ*~f�@��O��(��Uv]1��8!�Łӻ-�N�Q���f�}�R�>0��:��VҰ�{rE��%8�/H�-/5����v�E�I�D2�}�zl�Im��Ɂ.��,+���ɕQ����ռ�2t&p�/�ξiEB��7l�K��Ͽ�(	ÿ$��^No&��dq���W��8�W�<2�	5w�\�,a�%E&(��ܶ���[��;[Hj��Z��-!,,v��°�80��ޝ�g��К����(�OQ$�������3O�xm
V���n���D�T¨����` p.��|c��z꧁o�+h����`b3)v)�R�H� 6�S���J��/��+�-������bk�o��~s�ង��m��k���y+�X7��W��Q�BH��yη�oZ�{�J��16*m��G��l� 0��:ru�u�t#��A�9A~T�u�1�����{j4��2Wv��K�f�dZl�"�)����t=RN�؍����a9�cn�3q�x����1Ƙ���Gf�����3_�sY)����#�@6�ˤx��T (q ��e�����Q<���Ɉ��\�˓���S��M��g����k��0�}ԫ�e7�o\4"���К�p<����>U��� �<�iY��y4�`ĩ���;�k^�+-/.��3�z�������,��7��ի�h��ڹ�L�n�-�� �kf�%�@z-�b���Rƛ�>?�s��`�W~�n%�jEh�R�Ƨ��V7p�|JP+5X4������fx�|m8�_a�U�+���O���x
e�0!I2%qÉG�H�����-@`ʘ
�n�u������8T��[:��w$�|o,%@L7=�H�־�=W�e�Ԍ��a5�T?������s�kȝh��G��� ΋�������.2u��gއ��/g7�������v�T��ʫW�bW�<O���d�'ɏ)��� ��2��R�y�W�N<�\�g�9
Ե3���eJ.�]dL~��e�=j��gʹ���\T��I=�p�[���3hϞ�bp�_G��(�)M�g(G���0��D<Ih6$��Y����giH��pk$"�~�XE�j�ԫc7�I�)�1r���n��wJ���Ku�m>���|��]��j��I��)&��k�_��W�P1ccs���h�k:��+�}���&hh�*?)�M��br�wنT�=$\gk���`ӫ���v:��k1�&#K�_�W���qa><�֟ݑ�J���	
��X᢫��'� `������l��]���.�`R[ڭ�ʽ��ٍ�F���7ݧ >��B�383u	�,/�7�5H�J��gu�������a��7[F�vn��7�V��,}����ji�����_�gX1"��L�t��%=���[3���%+*����H��c�`ĺ�c9���XWj�¤���?��W���?���jZܷ٘�T�P���87����� �b9Z.���,���Y��jht}�ֳ�ʗB
}��&�{T�o�A(�eQ買��ù�M��)�I�:C��x6Њ`�1/��{��ZQ�JD\b)�~��C��_�,67����TL���G��,;��p�Ş�cN���aI�Q�� m&���(K:j��?�.����?������+ mcV5H�tG��?����P�^d�;Х�$($�$-��}Y�	K�[���(�����g�`���Y�	k���'�Ҽ$O��o䘚�YIZ��-��b�/ �����!騴�g��	 �x,�(�	O�a(�z�?��%��H�4^�I��)Gd�>)�*0�Dٜ{�[~���ߣ��"�_�?��D���e�a3��m�"��We|5ͶJa��J��w��.I��A�׼�Y�
��v	v����p֮u!5mA _@rbڦ��M[�z|��+)��Bk㰃�`0�*\C+nѣ��Q��>��˴1�X��K_6�2e���X5_��!m���}(=TF�]`yX�A�	��d��\V�Y4#h�R� ���G)u�{�-�U��I�h���$4��m̷2��.LY�R�*	�7tn�������a}B�fG,�I�2_�}��wW��{�)b�촏�e�J�C3:*�����ў�HJ�����T�
_%���)�q�06�=b_��F�Ger���0�e^��@Ȣφ�k���,Y���M�$�cD���tA�Y�*-�a=���ֹ�
-�#���&�5���K~���$m�B����p�*n�/��v,i�!{7�k9daJc�AwUڰU�R�8"�h��T���[�f�Οt�8�j���zغ��YF�}�H��%�Y��u
N�������h�`m.5y#��dbV��t|�;|l�E]^�u�	�+�3���A�#��f�;���9Z��'��[��]C����q���YM2���L� ˲0�'�������f��i���E����49�,G6E�2���� U�?N�r֚	Ѻw�����܁�r���{�W7��q�T�h���o��{O�K,���+p�$�m��)R}�4in�A���D�L�[&�O�_���XS�&4�!{�0O5][�4a�2P" ζ�H�~���Ml�	�����a���}�Ά��w�k"��yV��� V}]Nt_�+\'�7�o�4��}��qQ��
�b ����֢瑬Au�
<�䂜�<�~ϳ�]��G�V7]�9A:*�v⬤�I�'�oU�;!v�4�3�'y�r�f]�V���.��	���������m1S�Z�8E��C�ڼOe\�zC�r�0�?-(����jr�.*4+a$��O�"��͂u�B�i:?�}d�0|�7h���6��X5�����A�|x��t�1�����	{wO)��sx������ߑ"�f��.2���p�n�5��3	���]��]�}<
/i������k+�v��ER�b���5)�f]�����s�����$×��z���<�q���\��ߩw��l4�"��F/L�lN�$S����Z	p�Np~��w)%���ğ�����W����i�@C����{fՑ#=I�/U��U#^Q)V�����O��%J��@��ayI��T�4�˖d�s8�5��<�.�6���Ѽ���k�ޑ|6��&|�}��vI��AiͲ*,x:(>�o�"n9�A0n,����
=�`�H�?.;�"c����L�<���B]z��cP) �2+^%��%c#j9�?T���$�}E͉���ŵn�3�l�w>�غUuU�u\��/X��u+��/}�ԶĜ����G����S�1-��Ҩ�,���J8!����HNOFy\�d-��kI�8P�՞� 8֦a)LI.\�F���?�P��6>̯�m]���\��L�T/��E���1a=J6�~�n��0���y!���6s���N�HS񓊋����GC}�<�������7<��9z[�w��2F��*��7�\��#*Q#��b�P�Ɵ#�P�.9_4�*����f��?����2
 U����Jm�cR@�y
s܊7�����i�IJ�ib�8�ѵe�����x3vT�T�P���3,՝���E��h������ 6O��c�E܇�q�������d-c!���]�p%�2��,V� Ȁڦ����/���
��w�@�R1�l�5�@�]��� �{�P�g�Aݛ�bL=8�>�繑��6��NfD�6H�]�d@_�Hu%���
�����+��� �v;��F�k����b��%��ƹ�k����	�5��Q�9oy�Ľ����� �����`�έlф���+^Ly�|�Ê��؜T�1��(�����}���O��Z��5�Oeɺ
%��hA�!�-u��wI�z���i ��`L(����3�<���ijW�\���&D�,��8EwP����Mq'G�8���^9rޤ���mbf�#;��n�'Qˌ[���XAIP�r�
�Q~���VR��Y����
w� ��%i�5�V��؝���e��2�N�6�o�<��XS�wXx��}�d;+&Wh���u�-�3��
a�)HZ���{�׸PKL�]�`4�\������	�ŕ1���u�a�B]dusE���K��tp��X��{ڮL�@*�9�<����)z�a�L:_��1.�i����-����~�ٍ�������IO���cFI����#`�yt�Z2U;5�yD���P�M���>7���<5��p�Hc�_�p9���1�%>��c{3����0��qY|��l�����8��{ϲO�*� �V�����D�����5����Ҧ����a�Pז}��g�7u�J뺼Mэ�D��U��!�b�� M%X:.�ߐK�Ӈ���92���^ ��
[bv�&�&���Q����y���7R�N��(tj��hO�<���e�4,���H��EMݕ?�
�w��/)��#3�cw�>i����[�hm؅�-S��,7X���l��F}��X���R�+�_�gԻ�v�8���y�t�ޣ��D����^�/[*�d�_�g ]���nvi��m?�5���]CP�M�Zpq���R���K���X�-��	a�]�>�u��"����p�Vo�,���ٳ�-�*�������w��f?��w?�����A#�����xM�pt���G�e�8���9��ِ�(���u���9�]V	�':3.�w�*��MJ�ڐ�y�Z���St��U7&�'�>S��
��G.��&��$�E�ce�3lEGq�ăD��mdCJ�;@%���$�#�
B�\�d�ue�Վ��&K
��CN���*��tH�
����&�I�T�swz !=�ڰ7��U�{8 �\����Q����Ʒ����KY7G��
{���������,�E�FU{��W���Xy{O��fU�gsx��H��{�pWW_�r˰��dĭV�m[U�@M�[�R�xB��������q.��]��_�8�����%��>Ңn���|>����vY�CnU�n��ܐ��=ꏲ>��b7۸)4J��e4jWMo��ߔ�_dvأI�z�0��(���G wD+�WsK1\�4����#�\�������=��.���'�å��5n#[qR��9R����q�[��k�9�(}�mۺ&il��0��N�O
���i�G�p��A�=CxRY��l���n�a@ڰ��� �g�>�L�j��ߜet`J�iM��L�;.�`Ņ�~�97X��Sg~��.E�3`����!�P1�^)�qI�pw��Nm��<X�����/Sۜ{�"� f�}G�3�SL��-pK��夂��H�wS�8]�K�H;6���}8>$�1�j}�xޟgt��^,F�gi��n[��"�&��������F4�gMv�Z��M�(�̹:X���:h4�Dr!����z���ҝb��w������I�j��a��������m�j2&�S@	�}g�@V-2g�iM5�T�e�����VJ��%A�e¤Y;L�o-�`��Տ,1�n�k␛�{i��F��걔�I^]��Ip.ds!Aѳ�;�qd�WpO��5pe�������{}�VICouԗ�)�<2�r o�p����Pv!�,�L��T��ŠEXv?�n��r��; ���M3�6=+�!��<��#Z���9�pn�T��fǸ���"
�G12�Y�D��$�{_]Vru��C"�H*�gͶ~�L
3d=+0}P��Ȇu��󥘒�e�;���þo��T�e�輂|j�B����R�0����Gu��e�(u��[�"��� Cc�\�?��]<L<���>��bY1o���őo���tf�p(:��B��fLލԲg�J}����i����g11f�Q�m ���mj��NxWc�W�ࢻ�%�e�*��7P�t�F����Z���h�P*���@��Aw;ap�tPF�&	��RL3�������4a��=���u& ��8�"�9l*b�4N~N�Tk�Q.���F�Kz���m�a�_�����W�nQ�D3'�`�~����M�#%=$���Գa�^���&n�%[b�1$��wYW���4�Q�>�����LbW��"�0�(��=;��,��h@�K'��;m!a�d�hQ/jnZ@��i��5����z�9l;�[;uAV�3EB���$�2�~)}IJ/����1��M(-kc�VyU1�t�ʸ��(���
����7 L����-�,v�F�����<j;B T�C��5��0��yL$7����H��䧃�m��]�h�Z�����E��p����n�2l֭V�[7�4�N
:�����T�G� ����>iN]��s�~�!ipz
��"+(T�Ir��[r�u��3���Ϳ�#x��3'���o�Ѥn��<����4���?5�(weOE�T�.�W���W�<���
��PV�啐�X�p)P.�࠹ƄP�� �IL�;�S6j��\�Ѩ'S�j����w�i�7�����z,RnX��J����'ʌ�a;�����JڴT�����I2��$M�8ZgU�1?���sb�x�J�j"��tE�c=f�CS�Ӽj!�\�ȣ�9��p�h\$��/��8vb�o�Ϣ�z�0�=���5�+U9?��\Oe�V]f�<���GN�ǳ�*4����,���z���Y��GCx/�u��yz~���������h�� `)���}��7I�sT��#OL�%���QE'� n�2ؑ�S����.f�Ζv�{7h�\&r����my �-��d��d,h���i6�ք��?%�V�7�U@���ꕅ�x�P�	�{v�;Pa�`Q���Q�b^&����m�j���	��3�Eb�ߵ�yDC�.P������4���OU�n��mRpv�g�=Ji|�����-�ǔKy2 G�NVp����M��R:Y���R��\��*�r�I
lL�W!6�X:zL"�ƅ�ة_*[��d���e�_�az{=�o�ɣTZG䁜
����L�!�Be!� ��d��We�|��{\�:fC8C?��N9�9�"��.�l�����("��6׷�k9 ��zH����E��|���қ�m�U0�8��b	B�к��ƞ|_�Q����?V��FM�����l"g��%	�{�����o���v�Г��1���z�S��_oxO��,	AI",�����m�Bo��f,9�K�9���4��C�A��|�0�"$왦�!�ъ�y��ț����*��^,:���M���Ȃ:���0�Il'����W�<�+�����@������f�|G�D
��(���
:#�V����"�d&��e�2$��M5<k�_B�o'
�>֕�(Q�b�㭀<��r��0禢��8f�����|�N;CxiȨp��y�A���R�*kK=���|8�^^���{
��c�W��+P�����2@ci�OX/2=^'۰� �~e�U,gK�J��ɘ�#�J
�VXfk}�8X��RȦ��Z��@f����p~�ÿ��8�v�0��*3$ڟ������9��Q[p8��왈�">A��l&��,�� <07�������A����P�V��8���Nr�u+LT��H1��%K[�u��XZ�c��*���"�<I�߾X� nO7�$��
2��QX.7��^^����\�x�����($�-��9�eֆ�#Svh��a�rn����C�q ��W;�/,�c�G�i���o}o
:Xk�~4B φ����sOˑ�5��"핐,AAM��Ex��y��ݑ֠'���K>,.F��WL��ӻ|R#��V�C�<ߢ����U�@�>֑�ɺbE&�O�b��֙�� �� � L' �'$�x2~W��b���_g��u��E��TC�@Ƣ
e.U2B%h��]�PP�QΗrO���W��;�uL����?��>'�FG���m�ް�J."�m��ӾR�P!�!��𷗩FF.���3���&#\�9�����9���r4	�z��x�8��d�J��w[bߤ]�pՕ��2%�,�`�/,'����/ӟh���A\E��D'�3���|�=|5 �����Ё㳧�S��v���}���ㄊ�1lr_�x4��v�K��O��j�]�0K�8y�ex����/Z
�=H�@���ѹ2fG[%�Y��G�,tW��4���6�k�3^|T(�D�^)� �����)��	��"\b�I��L*�I�"�o��S�G�G�l[gTk7�C��=	�Qt��x�zݫ���1����-��
j��l�*�������t�b:������M��}�w
6��>!�K�LW0hi~�pץSI?���k��)���p�,`�� ~�9H�+c��*��@��,`�+��M��%�;�`�</ߖL�װ��7�.�� 3�Mehlo̪�k�S�'u)�����C@��E@������u5��6`�8��{�շ�����fd��y\����z
G��1g{:J�)�SP�`s��tP��fFS�<�ј�7Ѕ�W��	c`A���Sg#�~x#N�����Qh�^�s�l�(X@�h6`jG5�x�"݅����p��
��
��ؚ�,D�1��Nh|H��_��Q����|���!P۫��z<�V����9n�9z�oP���dDΓ
��N��X~�G����n�F���:}�N��xbP=���-�gߓgu�D_y�83G���W�c|�+�jĺ�=�<�hB�u��P���p۝@^-���[U��P�V�[��3H�F���~���A�.��&�x�	�~wQ5o��9�k���� d)���x)�yc%h�<'1G�!oUH֍��to����;2w�dl���`�NטeB�|}vڸ��ju�hJ��z��'��"���+�c�����託��/�������Q�{�>��r;�@��8����#�vw� {�h� TD��ƾf^��ҩ��zƽ���^e��Z}``��,2>1(��쫩
vi�ȝ���N�RH4NV�����熃��!^�K��F��(�SN���u�UjU]Yi^l�A�2,�#P�h{�g��H�_[K� L�����z��l�����6>�C'KS b�!���l~0p�β�JC9Xv��a14R%�oKbc&�jK������U���$mъ��d�J��$���Oe,u�;��
�&�Ale���٫'i��˽��p��:�?��j��KW�O
�.��[5�s
-n9U^�����*�z+�A�c�;���0���q<}r��1*0'+�9~{l��в?��ڥ�Ts%h����@4�)�^�%���fg2x���衰qFp��VϹw�_l@��3%������ �e�G\�T��΍��0 MV��"r�-�Zd�]4�-���nn�f밃��{�z�:|�T��#ݱ��v.g��~t�M��K���x3:��[VlY)'b���R��A��
q�y�wC(iC�,��T������TW-�o�?�gJ��	������!SB��f����	&3�V_�cc���@)�$a9k�oT4�����.Y�'�������CѴQI�妟ȭS_���P�2�b3*�١Q'{����%l�,Z��6�T| ��]ؖ)��<��KS�=ER��G�P�Q�c�hP���/7��G�fˇ}��^v=���y�����d~��SJ_�Kt뀼���^�EFT�t=eikS�A��֤wo�w�;�\g�M�)�ŭC���}�V��G ѢB�=��F�@Ub�%w2�	�=<a�����o�6�~��G&���m9D���X|b���86^���J�A��4��:J	��+{%��ݶ��l�����6h�e*d@q]T�Y���]X���
^��\Ik!ʘE���5�?{X,���&Z�7����ƞ�^��E���[�ߥ�z�t6�#�spO��ʡL!�XĤ#H�품Е ��p��/p�V
� 1��2ʑ�#]���^Z=k��W�2��֕��u&��I$&o�h�ܱ"�+ }���\�4��q�T ��t�G.`v��N�{
�Jĩg��1A���^�<ހ,+b��m�[������s�zF���Z�m��n�X�[�D�����X���fMyr�K阾�V�	�O�u*�ab�&i���k����cZ�����������ڝ��hu�nzh����K�v*���54{{^6�2���\9�٩��L=��TNT��5��PXi�M>����=(��e�Ѝ����.E^](��V�`$�s��O�y`��Ց�l��m����U�n��!=�϶��j-�<���	�����FW�[W�/5�:ə�J����6��}�/��@�5���𳃔��q�e�V�@F�ѡ"�U!~�[`� 7����TbI���7d<d4Y��}�b�.g̺�#�jZ�:x[-�#��3�DK���.]��H�5+�ꦸ>%T�d����D����FLˉ�󉙐�Ƹ�;�[o��\���epY�$I5�_<"�a�v]S��fa�W���?d��m��31#H�]��0�fN�ͺ��^�I	��������]��W��S�g�JFd�b�ƭ,w��s~G�bl�HL�H�fN�%���O[e_���^�)�4+��F���g�LY!��8R�=Q>(���)��u$���`�Vb��#7D�v\�1ʲӌ��2{���,zu9���=�g0�AI���*�߳����w��'>r�-}�)ǇС�������sa�����y�'
�w�fy�J�5@0��������#����������ǣ��䘭W��#�(�{�x��i5VB �V�����[�+ R�FK�� ����r*�Q����L�H�[��?�gc�w�2�� ��蠒���x�;�P�K��i���	.����4��i�g���?��s�qmN��*��mQ���-�"&dM��#�; y�:�p:�_L�����\�sV��-B�f�88^���{k�����IE�Ee�S��̒����*�Wt�o� ���Oy���,�@(m�NT1�[���+�ے�G7M�O��h�	�/� p���A������k�Fw�[��_��^���L!NH��I��]n��S5��xv�PpM=vΗ� (�q����oJp�Z� ��k�=@,�Is�2��oP<�ZTآa���>��s!�%A���@ҳ�?���C~�����E��<c��8,g��+�T}qv�\k�z��(�=��02��*��>E���s)H���y��v%��W[]�ٟ_��B0�{O�F"�n%��l��9�>���c";
����й%��M2�������� ���* �ʎ��t��}|	U4������V������]g\e�fsQ��Z=kV�Ag�xNmi�*��>׋������q��*~<4�ߪ�p>\Tmv�iA���z�G�p5�ʊF�mvL�6W9p�S�5P	��-5���
cB\��#r����Bzg�'W�Z��'íG�s��lfL�q������z�5��YS+�3�r�ˇ�*������j>�YJ���RH�f�9mf��"�ngߩ���(�@NV��z�?�vY��<1�`V�h�=�%�h9Mj,
�_Sb����z�C��Ȃ��[l��~�>�!V���d�n���)���o�Tg�5Ԝ���yS�	<pH�=���,�9�D��%z��U�B�a�z�҃�K�LOG������%��;����B��%�)�)Rz;�<����^�*!�Yuȭ��ɻ��0�X�#t�6)=�U����Ӵjܩ�cS�Ck��Eؐ�><}����6H�\�6D�g�I�vS��خ�/1�=�f�[̲Z�C�m/f�:���,[Ĭ}߽W���$@�u�Öx�}�>�4��TA?��9���v�[�%I3ꨃRuY�`n?$o�w�ܖnR�e�A�!�Uo{*6�*�:~�Z`�0��@�1X��t�P�^�VD<��ʝ_�B6y�@-���n�/�����V��d�3�B��9�=l!W$S�V����f�v��| x"�܉	�%k�8�,[�jm,ۆ���Yl>:���D�ؘ-�M�YӡQ�cҥ7�w^�Ip"~'b�͒a�QI&���+����T�c�#���^R /m��K�h.FSzZv p��29Y2+�C��]E%мKU)�H�UnE�~Y����վ �b���:=C����bũ`���T���rP
:p��=d�(n���e����%�,��<h�rT�ފ�UM���\��4��`�N�cD�@�,��߃%�B�jY37��|�C3�p�נկ�\���s(^�!1K{�C�g��L�_�!���&����Zc\����#�߶����v��Zv�W���`F˕Y'���=�`�0`8':���ҵM,(O3�=/M$8�������b6����R�~�_�>u�m�m�G�!а&��%יu�1Z ���W�����~�*!���n��&�j�3���IHS>����-�����v�2F+o�V����%!J���C��<P�jw���2��۽E0�sB^;�˗��h�������K�=Ԉ �j7z�����r���@�t�H�S�Hn+D�M�I�jT�.�-�ל֭h��ވ�unʁ�T5�x]����lh����$�l�*�N�Qt��+�|3��?E�Z4��tK�dyn�4z�ip�>��@���B�WH=�[v�q�/a8�¡_E��ߤ0��P����T���n��I���d�]�¦�M\
��͍�w�qmr�'�p9��?��|q"W���5D�r\2�x�� 5����?gD�A�~�I�+�4��=�N���Xќ���\O�R�}!�_��ڛ^��aA�NS@Ìggֲ��ohZ��XrV�8�"���B��=�T'W�+K��I�%[a�"�Lj�dX��u��h..���0�:2��Fon sۓQ�]�hc���]%�6I�F0��	&<�V�^`@��}]�XY�(����� ���e�PaAe��(uCD��P��������r�g���"��ղ"1:O06�Xw0���=�� J`�О'����Z�� XU�R~D�3�)
1Le�}i`����ql)mM�%�,��ӳ�������勣�-#�y�Q� �;���@Ʌ�B`�C����E���-w�Bg.s�?�|͓ڭ�J�*�Z�4�o��eufy�-�����<���1�@n�T��U��b�Z{�t���'��ړGTR�YF�Њ?R���ƃ VY���V垩�48pQ�ny&�B���B��v�ü[�O�6��o��[v�ٳFj�ZÃk=3ѩ��nl~��)���I����
bh���N�3M��FH���<
V]��=+_�Dg�o-_�?_%�- ��x����O��e�Ex싸Oo�DH���\�TX�W �dT^�S9ٌ+[`�D�u�r�s�7��v�Tnc�>�K+(���ǘ_kw�}ܧ._���1��pW`�퀜|�䄻+��l���=ǈI�<��~���i�o0��c��2
�(�c��C��1�p
O�-1H�(�L	���r���У�\��:�'���A�_`7T
��x(
��2鉂���{+\�~2�P�t�~'�JW��������\'4�+�t0m�1����0h߿��@+q�� t�$	�%`ЙRA!=�^;X	!,#Y�,�X��85>sE�I�>§5A ��C��|3a�m)S6�z�:���Р�BV�������aP�ڏ���UB�{=-�`���#ל[7���'Y���#��>�HW�+��9�� &�1\n���k�aeq����D������u��mm�)��꬗o�v��B�x�alkI���z��q&���l��(Rش%� z3#���l��;�4����R�	��:w1��|���0�Q��9o�߫�3�1O�)_a��9�]��e@�7�2�>_V�� I̮4������-�e�Ν�.�-��_14�#ધ���˱�������:���v��QM����i�輍C�Bi ��3*Yf��!��-�+P��VD�%���p��y/�*4�g2���ອ�4\�(���k��}��R�
J*c�P�qK���1��5�р�H�u'�Q_r��D�,x�[\��]�\5�<���o��&�=�Fv���ч{���*	s���,��zn#!gB�=3�d ��e��G�ǷM��3���V���&D�\����餏��
#��.�0��z>��s7�b{E����Z��F�^F��`�����:�G��6���(;�c�v�:����EY$��E_3y�8��ܜ����
�y쭺��hǼ� d뽄T��Bj-��1lX(��:Q;�����[%&��W҄�k3��]�������kgtOAU�F��X!t���*���vF�p!h�y�-Z ���5��7�==~3�{��x'	ٱO	{�D4��fD�������;�j�%	!n�X�n��m|��s�����E����3O0P�6t��`8�N����;�5���jSԪ[q�?Vj��~��w���%Q����>���:|�U����{2�H�R��Z�t��%�����;�fX��ro��4�sw� 0z
I��/�٣����1���WP�`p�C���{�o�2��IF��4�]��>�vj���x�!��ݙ6���Wޖ��D^����0��cQ���F۶��f�va�b7~�3ݵ?��m\L� �b`��I�4�,d��guh�#4�^k�GUr���#���ݳVC9>ܧ�S���D�Z�f!���52�Y���7��|�@#�?x�Mpz�-�P�H�l�~݃컆S6�A���/���P�"��>?2�e� �%���uG�^�}ٻ���9 d����qO�d���ɯ�6��Q1-U�ℭ���:�ظT���?��L����J�/��z��#�>��	��d�>LY���A�|0�U�}qL׆M�Z��f�N�\����])���5��]���F�p��w��o�r�lqs�ћ��_�L��~i��g������?i�C+�;���܁mE��h�(� |�4�Y�J)CA�@Ԛ�͑�2d�&|Z5�H߼k�E�*Z�����{m*���iYu���'D����>����K��=f����]D5[�U�[�+�1L�w_��0�3�%��Ւa��W�A��P�Se۫��U�2�cJ��F�Vơg��)2꾃�4�7���y��-��DS��s-A�
�̐7������]g��Gap�~#b;%-S�����e����{$����q�@E.���l�?k.OP;P��p(�ѯ�w�J	����ӫneD����}�mM���?�@�p�3�?
.��`Cx7ͦld�R�l:�$��W$���I�L�t/�G�8�2w���v:ѫ�/�:J.I�&G�=$�Z�m��M�0*iw"��3�L��,��J@֊|,��{׮�1�%YН0�k��^�ζ�;!��}LzbC�D@��̜/x���Я3�?yu6��cBኴK��B_Ѕ�؟�y�U����wRjV<���ƅ�9��_qV
mA���t�G���J��aP���l��AJYՊSi`Z� ?C#ZR�a� ���P�a� $i������U~�ƐT��J��6
V|g����4��J�ő�B��U�KD�+{Ǚf�5����c�0Q��Dy�LQ �bx!j�z�tS$���I��0�0Ѷ{]��"��f_��?ڍ������u�Z��<�7��rX����Y[I kq2[K��\򅶢�#��z#�E��
l���;�<=�?���N�G�g�z�W�����/�(A�'��j�f��b	�FY�~^{BCE`��O͍�F2�y���g��R�_X����*�a*
c';G�G�"�1���"�!`X�uAiG�a3�v>*�aO*��o�[��YE:o�w?��oc�[�{�����(F��fM�T�d��~H����P�/�BuyDu�g��M@�[jB �j�p� ���Y���Px�8h@��<�q��T����_�b�663��ƻ���^x_�����A���{�f�vҲ=b��Z��<FgT,�����W�o��9(�z�_x��c�|(���p�C�l�-j�@Č��n����b�(9Y��(ˣQܛ����~pVum�L F�M�� ��Y=t�3uOȼ����R�]]8ɡt��+�t��ɳ���/(�x]�;�oN�k��3��8뙎FJ԰k�#�b&b�:�)� �n#�'�>�R� ���(��E�u"�h8i���t��Q��SM?�u��u�1/ɵ݉��mR�����0	~��Rl�V������D\��N&{�Ee���l�Т1���0���|���¡q��/��'��d���d~��'za�%cVQX�^�� �- +�_�!&��'���c|��5�+J>`�|�R�H&�@��&��� (��I��P�)O��b\�]�
l�|*���ژ �r����E.yi�m���G7󨧓iu$�,�O4��"����p���='�-�i����#��$��)���Q���H����>eօ�E�km�JOϼ��l�ӢzD_��u���*W �r��ώ���?[D�Z�6�Pł����M�á\i�#��*y1a�a�`[�(���lӧ��"�E�Y1��_�#�3]�'��V�pE�v)zG�=ҝ]�<�7c���r]
�����9g��9������ jƧ�W��lN��MO�sRQ�frٚ8��b�^���˾� ����u?e5��Vc�M��cѡ'����|�WI�5S��UT�ȝ���=-�5m���#���3���}T�\>ne��D����F���~#���U��G�GL��)�l����0j��+_�/ƺ�=(A�W�EO-BC�K"�		��ʯ��� <<��j�&��R����k5�b4hzD��y�`n�S!�D��䪃�: �}$�<3�0�1��%���6ڄQb�(v��uVv�ӯ|n^��w/�q�/Ro�/�T俗�r��~�N��� "x�\��E���P�8t^�Zѯ���No��?�_�a�T^ה���b���e[nw�� >�����*|ZD��Ex�ls��~�Q�&�n��E�3�G�]� �����@��ޣ���O���1Z�*,�����yN�?U����Ǖ�����T�"f�m3��;i;x�|��X�������yD�)��v��Lmi�Ϙ�`s�K������J>q��"���gÜ;Z�����d�*~�b����:U���E?`i���ˣ�@� �0ip�C����c�QԔ����\R����t���{>�⩄��S-_Pw/��R���􌍡���9Jt�!\a��g��OG��Z9��X)���Q�*���k�:<HD�#���J���ڏ����q������d��v�e��������T)cp�R�h�]7�$"�i�v;�5=J�x3q�ea?g|�|)�e�Ņ�S���7�,����PS�;�[X�N�s>�G��8�$��T����0�G��hϤ>�,X�m���6I՗�e�%�;n����/#� �h�8V3i�݄>+CIYa�FG<c70W;y�5`_]0$�.�$�x�g 2:A��]�{�Wj�Tv�	�ؑ2z~�8Ul����Š��#�t�VP��Ƕ�~6&]���xL��XBz�����LI��s��B��IG��� w�D�S���ūhf���_uc��4t~lb�4�YYi�t�?:�5�u�]��4��G�h*�?n +<�X��ג��:����}[�:�!�\=��:K�pz���� �Z�`��EHh��(Y��FIM��sz���?W 8�+�lx��l���=�S�[�+�������&b|�^Sq��(3W��Өb�a����zW}J�x",�	�$6���zS ��>�6M�1�=��Xu�хa��h��o�+���d藫��6B�V��,ɋ��7��˟���8�iE[��ӧe�d%���rW��9�U����$��D��m�FR�rɽ��:"���Cx*]�m���S�|0n�dF��"���x��H����r9�_��s�8��y_��ͫ�ۊW|�m��-o��n�$�>�ʏzx��(
B��k[E%��/�=����/��}�ˉ�E�LQ��r�8��_~�
.�H����o��;��tz^G��>Y��d��p�8��jlm$^�����XD�0���c��8���./�����Gmپ�c��t��x�V�Ll�z1�9EݮV|C�=����8��h���6_���x��5?�J=�Ƥ��3F�7���$���G�0�P+h��T x�q��6�,ju�0�H�� �"ֹ)ʲ#tN<*��N�r�H��Lz{�U��9*�w�uE�_��:
%l���`X+NZ�;�,4��fA&��7ʂ������b��Y�}� �g>W5Ӓ��zX6J���wT�x���l�x�-�'�:�W�J�ir��{�����vzǵA��BSo����N���%.?���-F�"b;���������l���%�'%�x`ڑ�6C+�e��ctD\�%B��Xa�@똡��[� ���t5�B�!C!�9��ã���#���c�@����;�l���q�� ��ff����wt,/u@<�._������n߳0e����ޘ�x���kt����X�hl���L�j�a���v3o�C����	���V��L�@��!��CU�|���{4� �d�b�@��~%�/��<u���܁L�1�уX�`�w;6p1t�ĞS�ח?��K��m�>q��eNP�zWc�(���	�o�-i�W�4��\�&�X%z<l�#haFW�����ؐ�<ٜlM( �� ��(_��[ɔ$q�y�I�g����K�}ہ�F1N7���U�eo�Oåq�Mo��vө��UDy��K�e��E`	n�TKfx��`r��X����+1�m-CD&Z'9Cحt�byVqVf@ऱ��e�f��+@P?�ӭXX��=Fo��%�D\����]��A4X��9�!�3b�`��˅�:���CZ�J%	[��_�Q�J��*�@7��'�8�w?�X��C���&J����(���js�p��*��o�kue�~��d��B��H�gO �t=[콞^��-�H@مnS�����C�.H(6�=iB4��O�X8�B*N9:4�X�F޲v5�WS�y�!J�=~ ��BA�g�땘��:js嫛�����c��A���e&�<%M^]�3?�kR���Az�Y*�1~oD�P�%2u<�^5�&���6�����瀾Ѭ�+)m��*�m����^-yA��۲�W��� �����8
s�U�diƂF>R�ꩅ@?�M���]��V��N��z	�+?�k���X��l�a2�C5�;0�Q�Is��-�>֏��UlY+�e:��H��]�R]����)�$	H�IK_�!P�ZdF+�2��5Z��|h�v�E�0�G�Q��R�y�<�u��[)nY����5�i��&�k�ҍ���z�1%���K������ɸ��h?3���R���vt)D4V9N('.���9*N��o�8(H��UOI��a�����	�P*ᒵh�;P���,����S笏����#3'��Qv���qr �ޖ3���y��DɊn�B0����M2��� �:KO����[z�̕�$�6�h��H�b��䶪9n�Bج��g�ݾY|�df͙r��3���6�q�5�9���G܊F��ԝk�J
�z27�;�', �y����ݻlڨk��#�p����i�����#{E,1땣�?��}�8�;�H-ʔ��^All��������l�	$&�d�⃓��d{�(�!����B��U}!�ǂHdW�V\:�抻�{*Q�\������#`�c�����<�#N]q�^� ��ERM��k����C�� �S�M~'��ѳ��0rN�P�C,�*��m���w�М�q�ւ����J}�E�ؘ���>��Z��oq�61xa�DQ�S��m�P)��	���aM1��S�<d��{�_��?J�OYy����@tS&}	����t٧2���O�T'�jh�8�6¨.��XЬ$<�ܥ�n�jC2����A%��~�K��PΑsA���[�s8ץ[6\UT��}�ʡ��n�F�$N~k62[J�����&'%�R���Dk�:E����"��@��:�q�Po�`���R.Â-W9��@�~���_�4�_Ia��>�����"���>9�[?'Ձ�$!K>�<�!�TB�Ǝ�����_@�^��>�*V�ēg�7�A e{!r�ټC��@_x���^���qJH_)Ť6��I�����ZGXѹwy]��r����~�L3z!���F��6H!\�(E�z5��Ǭ����x��> ��ߥ����O�+�tZ�U��Q������Up���U���N[�[�/ik����Gd,@�����Q�s�R���Z�5dϑ����L�L#�z�Wҹ�5��1�j���W����Y�� c���l���W<ppC5X�)���bp����G�$Z�bܖc���ʓ/����|U	I6<ղ�� v�J�o^�m�3��������P�%�����) ������X�A��[$K1١��'Ӷ�ecN&��)�$���{�/����i/HK�r������UCghK�P��,�r���%Q
�p���[v1-�gBE��a{I��`�@���p0���9���� ��|s�V�n 6�g��5��Ńr�g�_~I�/��ht��'k<B�Z�0�k���k/ ��/b�f�n���c)�M��M�`M�Ȑ��(A��Ξ�j�*M�AI�L�:ZY�{�dl?�*(T0�Jh��%��0}YD5.!����z�2:�NAȹً�5�ކhq*=Kg�3�d�we4A�b�(����^.�����5������}e��s|%�?�lv(�l�����UEp9��Uz�/�����S��o��H���~}����9"�U�u~|�r��6r����.Y�$��	ok�p!��Ml6R4(3B��H��������Q�z1�&E� U����,y<S  I��竊P>دsS�<b6��w�<
���Z�z�
'�Ҫe}��]!�t?�Q��񇃪߼ٸf��dav���[��
��iun������s1��_/H���X϶�]wH7�W���}H�|!�:���,���U�h#�+n.��Re	�h�?���
�P��;n�id�6‐��η��"�?X�\�G�7�O�,\~���L��ePg��CqO��8Ì�`]=�0njm��.OIb�|��gm0H�}�HnO��3�/�W��D��Z����9����S�530�$��;i�w����b�0Dz+����ӻ��pv�Rl����1d{+F��D�'hDE�R��~�N�.7��$nx7U�����>#`��E��9'���Xj���}��ߒ䰛��p��q���åb�~�?|�ܤ�����4[L �W�S:"�>Rt'G�,�T\�����`�H7#�b��yz�O��.��\A���G���5�i?'�[~e�K�b��淈��J?��DW�ʎ���S�v �����% ���������	^K��Yj<���Z�$qp0o�|���B�?OM��a�ȪN51���Oa뀵�ƹ�S�$ڕ.��7����.ҫ�xo}H/~��b�Y������8Gĩ�5��;"������q)MU�����}`��!�-����V��mR���A�_d��0P#^Z`q�c[23����G�����N�5o��/�Ȟ.�u_�j'S4V�Ci�x�;�ҠuF�|`�q�k�t����������R?Y^	&�4N8,%�ג��
my7ߣ^��]�e��`���.v8�ub\iߝ� ��~���y��s4o{.��\C�˘�=���؟L(��_ddE�Jʦ$����9��g��R��&��a,C������ܛ]�ؼ��M�&ܗ� y1?`�?Ԙ�Hy$p�\Ĭ�D؃�I�%�0W�|ޫ��&��U�xkRj{!�EXY�7�����B˳��������g�����u��%"I
�y/��x�,���������m?��=Y{��*�7[ѿ�z����,��.t�v��KL���w�fJ�=O��`tUI�K���<3��u�PuW��*l$��m�:,I+���O�>`v0�`Mh�l�1��g�x�I�<�vT�1�F�;̠��QH�X�{N��^��r�|��7�;� ^,CQ�O�_4�5��?`Mآ�-诱+hs|�S�T7ӒR�Da�ɘ_PArɋt��I��MxiS(�Ϻ�Ew���'Qb6���Х�9���:���K�Wx�R��T��cٲ��ƸǓ��ג�A��@�Zަt"�pLs'�揽�m���b[���e�wriA3�e6y�6�u>�:/�s?3���I���?{�z#�1�i�*�zw;MG�ײb�$3�C��܂zJ]e��������IQF|�^ʫ�����f�=}��8'i���@��S�X�F>Y��e�Y�%X��y����ݓ��娈��s�V������p���vr��5�0�S}h��S�~s�>yWC9J��O�$��J�1���FɃ���mK�'`������G#��_�������;m1Z�(��'Y�6z-�}%�8G�'���`o3�}ԋ �1 �H˫]�~Η�^K�Mx6l��q�S�����v����5���|��͋�k��&������y������P�\���B���J����U�v�E�>(�t�tZ�
!�g8��'O��&d���p���(r��@�W���m��X����b�̸ˮ��i��p �\)�r��K�b�ģ�OQE_t������-��Gg��~�#e/��gH�W��ː���Q���A�K�!�|��`k��d֛l���#�fJ^Q*rN��~5 	@�y�r	j		��>�0O;p�d��x�)1l(�Ym4r#�����U�E�,	�T?�Ao�nj<;�� �v��C�j���l](��><��_�#�\���c��*Am� �C!)�z=�&�T�ǎ��v��mAA�e�Q��߸Iӈ�
� Ft���L ȷ@y�֊�v���AF��<h��fUI⼉��2��VtV�lp�m�$N��>k}Bz$�F�`������4��w��!�Y�$c��LW�VN�ŐY�{|O;��s�6�����>c��Q����ԋ�t�#^�\8{�5��u�d
CW�ʦ� ��{Yl:EMD��v`�6��O�77���E�[��t	���d���~�w͗�����,42@<�z��0.�s����J(gI˪�n�Q%��wg�,���={OB�"���5t��2�aZK�;J<SЂψ��*���� �cX�%a1]�WA��p�Zڃ����XY3���1�+�3�_�{H�V<�~�l&�v�Q[y/%G�U\����o�K2JW����R�'Z0圠��Y�_RҌ�k�� z�5S��T�ǱG6�(�r �*�}E
z�l�]?ϑ����tb,y���,����Ι3��]�$��Oߏ5��<q��%T��2�H�j�(��؟ᶒ��;���U2�'�w��i��J=���܊a@����y���)l�������a�t&��s�z�>�W�����QK��`a��͞�ܚ�Tn���,*iR�m7�4N�$�ӚV3�����/�N#��J�M+R���i�rV�{tyH��ѕ�cN�.s�n����Lw����1Lf㊣��LL���@�i�Ku;D�Ӂ&���۰��^lƓ��r?&xU�A���D�݌�Hր���Y���OJ��Y�r���Y���!����������~`��}39wx �ʓldƓ9Ir�����X�ٯh�F�TP+F�L�b�� �O@M�9Y�i&���+�X<[�\J�� Z�L70�y���R�˞*����&�R��|�\V	�Ñd؈D�~�W��FL� ����І�!���x�5?q��u�t�iH/�C݂�6N�P�mg���%�5柩c�?*�Cv�ZX�e���vǣV��F��ż��Q���`�=��lY0'�=���&�ԋ^J��^}��vg��bJ�d�c���a��mL�Zm�,P���C#�L'�/�*����>z����S�Z�tq���g;}0R
�����x��[JW�����n�����LϹz��!����.�`�"�dx�>����f��RO1+��x�O�lG�h��ԉ^�..3R��<��:��XP�V�s���]4ױ�*N���*&T��ܧ|�0�-C�9��s�S�޼�Dt��I$4��JR�cq�J�;�V�����\	�v��˧h�!��ت瘐��q��p�PH�0uE�(:����l2���i��$�oT���y5�~@t3��e5C��iT����C���r�R����(���ߧx邖�3����	|R_xM�4���a�I�^zQ4b�
��
]V�1�����L+m��.,����ulh.�31�HX�$��S��e+�a�mP��������P!o�Jy~�J��N������5��T�V���)�B0͑ae�g����f�}���u��]3����B^ӈs(�Q�l#�,�4���ry/NO��a��<�3���,1 ���0��>�ľ�hH<@|���@��ڴ	�� �H�u�{ �Z�FP%K �}	����H�Nk̎Gƒ��Q��xg����iV՝d`YwH����t��$Żj�t\�ょ5A�q�7]G(/G.mf��LN;��ۍ`y?�i�7'��(d��v-��6�N]�.�}C��6�X��[�}�ev�����9���G~��}����4>wn N�2�*�v�����m��U5��b����2��`	r���S�Q�鳳�]\��J�yN����RH� �Y�K b�<��6&p#3�kB��b�v�x!��y��r�o��sD�
y6<}jl:s����T����3i F+næ�కңJ�؆ɛ�t�VIa�E�2�G��P�y�}\�bSz&nr#�";� �`�92+�c4�K�Bc� �����].H��)�rQ'�׻�,�)�H�S5y�)�������t�qi#���9�M�O��B��ڲ�s�D��;���X�S�C�X7^4]�,aڞ�jO�ʪV�[�!����4W3?Óp
|P&�%�}	T"�*���mI��>D�/���=�jJ�G�y����k���srD�y�����
Ռw-!����W�Y�7�D�*>��,��a/���;��7�s���*�^�;�o�vz(R ���3(����H��&������������J�>'���Dm^�<���X��?���s�% .YL�`ش�-�6�s$�i)K�C}��F��3���aW�{��5f���`Ͽ���<��&�D47�\{m�P��˸��8R:�85�'K��Ɋ&6��\Am��,1������q�Ea��@5u�8=tc�s�4v}\ӄ�M�5����#��?i�k4"�kT�����R:�5�M�$�.7"�hO�
c=P��	c�PU�s��q�鄌~W��P{?��w�Ew�v��:l����!��XƁ���T���I��)�#�z��I�	
	�pq,*�dAa���e!����\Ra��QM=F��m:=�9�U@���ڸB���1�L����*A�N��v�φ����NKs�$���sw��6i�$y%x,�k!{�]�y��O/Ҧ����˘ ���\�rUe�S��{-@���x�w�'�Q,}G�y|j����p��.S��؃��pɷ�o�q�.y�<)��V��W8D	p=@�2�y
xī0���2���A��o<U�G�G�S�k�,�i]?g���_A����sG��?g����rА��i(f�^�	��������x���Vŕ�Å��X
ڡ'�"ޤe�� !p�e�N}�!�A�=C�����i?߼fe�Ѯ�^�V/*��"�2����0t��0�,w)�j�jb���a����U���-H%F�T&�<pH,X��#)����2��H�e��G��!`�9
x_]qe����n.�[�"�eh�!��9��W)�l((��@���C�?XQ�y=��P.U<��_�%�{C���lh%���&�И���*Rƾ;���S��ıĝ�Z�Qo�!�3,3�[�
O�V�T}t+	�)UM�ˬ���~�QXsfI��!I~����!K����	����,�	����UUQ+�iń�o�w����<�2Sb�Wb�54Z��m����
�P�CWh_�H��4i� �jH�b�F�+��JF �:�^��b�TK��N������U�w�������7$E}Kyn��7�ֽKrT�]{����-�TM#"$=vOy{fp�fQ��e+�Wy`�H�o�G�i�*�K.¯�� �}8/7C]y�S��3�A-1�B���o��3����� A`�{Ӈ�}B�VoBQe�+稪Y9�b��(���BP��F.8�4�7E�:�$���րn�V��[`�/^���AϜz)4�0n�Y~��|V��*��/��I� wI�U�	�;Y�ct�6_�(��9�ʹ���r�!�ĝ�E�C�a�tҡ�.�h	B�'5T��B8�}�#�g�Z}��;��_ԇ���e����P!nE���Sd5k�Et�����i�Q�L��Ļ���|���G��)�)92�r�u�g��
ESpĐ�Gu������o�n�`ܨ�t�� o�%?饐7�����$��rA�0L��Nð�z?����bcAstv&��\Th<��}ܭ݊a�Z�ښC>���)�'�!LeȠZ�ӵ������L�����BeXߛI�7�q'�8+�}x�����&��ت}��nK��OX�)�;��U]0V��./��oL*c�&@�x��MzH|
5ۢD
v��ؒ
j�I�U�����@��}�JtJz�/��b���'�/�`vQ?�ߓ��t�e�8*0��y/��g4��+�q��=s��{�;@+W��k(9D��b�O���ɘ���B-�'�13=���d</[�1�qA������A���7)��� p� �VoL��$.�&��LJy������d<%���s���V\�(\9R?d�G���iL�
��������	�dp�O��Qkٳ_�
f�h��L��M]�T�^Q~��xU
i�쿳P`�����i�xe����3��US���HQ AҮ�)��zT9��6.���Z���<���~tF��g�΁�8����m�0z�J/��̤Q�n�i��J�"�>+���@�R}Ѩ��c�{��t~ܛ�";JS6��&rT~%1!l.86 QX��J��JJ)���z~�z����^���p���o��@��d��g��Z�̭u,e���]��i��,��K�^F�qC1�Bt<g[��:z��z+#����S�fRr��M�Q�
��^'��!�m~���6	��t��_as��F!�y6��.&�,����Wwٍ?^��B�4ɋ��G���&�\!V 5��}�ĶL�@����!-�o�62i1��`�\`±�͛��.���EeH��`c��33����_j��F�������4�ݏ���ǔ�v����6~�3�@�ʳl��~�1S�I��(]ݶ�+f�[���41ƭ�O�~�}�v%�~���e'���r��{�,Z0)H�����F�����J��SSU�T٩c'�$�2��z>I�$b��/k���OB����>��zA��]���n�t��#�##'R���v��w@'>c�|�Pf�&�`�8����/�c���S��N������;�C����t=�y�	3و�Q�I�aF9�^	���Y��- ��_���b���qf�^�2��1i�A��ją�B�����߲ϦNw�̷b�8��΍8i��^�(ȃ0�{�B�l
��}��V��+Vk/* ZaY��4Ni��0|�]Ց>���*Q�S5��1�GqM��|�l�鉣{�0<����rFbJbR����D���f� ���e�����x㙎�)<��U��WΖp�R��Oa^
�lϡ惡�e#_��.ǱcI=�l9��g$8��$T�Y:����.s{<s�%:*i��"tC��-z=/ Yk��:���]Ay�.�\���2�2��`����~8��ˈ\nOa�|���7���w��o�ht���Unq8���� �a�f�K
zA.��B����FlR�o��M���`	v~Xo��{Ni�ġG�Kc�2���$Kv�����^�ssp���c�:z\"�ƴf��|cPl���g��G ����"�)3��B=By,-�U5�L���:XVG?:]po/*���iv
��*�Y'0-�YL��7�fW���u�W��y�v��{q�e��c�I
�+phW�v1qm\�w�@��7Ӱ�'d j��}ԓ�KU��ʾ岷  lw�u����s`Q�.B�J�����s�`V�����R{���ۏS�ڎ(��c=d1��������̸�f�.��sk�����������#D��G)9���r@(�!e&��,�������c�LSڽA��������T��R�yc���#�@!��zyMjo�� }e2��5���m�ُx#�Mq1M2J�Z��,&[=�]J�w�n�#x?����"|�'/���&����h�6�&e�C^�|�r*p�!;�'M:�����>��\�{w_K^�p�)B����7���ڨf&!k�U�d�q��t�s�KV�=[/��4�&
0#�u�ä��t��gp� =vB�2�m٬Ǘs���X�㞏vZ�aN]�Q��qqv�������v�k��;�W�+(�U�'����Nԝ<�	�QB���PQ�\�uǾ�$]֬��n���j/a�K�݉�����ݍ��'Bw������幝
g�s�D�P�B(i���nM��qN�)��w�S��mO�h�GŅo�o���1�.�	*B#���`�3��f�-�N!W�.ԭ�"u*���eBq�谊�n�,?�~8��;��$�S�����0�0��5h��T#ٸi@�3����A����<�#A|�9���g�v��GӦ��lۆ䬔Bw��Ԕ]�� �v��0���t$�A;�6}�o��<�q�4oʜ�-�/s����E��"d�Yha��T����fZi� �W�%�����쏓U
��6Uy+�ag0N�	���v��J��. {4}�N6�6�0;��-�N�1q󢀤Ѳ�'��z�W�����,Y�+7��5s��%�����c������B�<"���ye�2���4ɰxC���ZL̹�jJSЌ���������no�,<�k�� ��a�nU1{Z�䝘�<3\5����:>-'����J���E�K%k�?|��=����l� d���D|�%�� F�"��[�)�*csHfw�`N�S9����aS�@��R6�i�g$��ѨV/��ԇ��e�<h1[��3�|?^���F��M�����4߸2�B�z�98��*y�������{����R�9t�q�=��T,�	(�R�S �Q�f�5����P������;7���΋�;0�t�\e�auւ���6�&0sc�޸J�eB�ubO@��-/�����焨���IW3h*���+�J1���";�d`Y�x����i��������Ѯ?���k���׷��q�ԑ�E��u)�w�1��%�	s[�����e@����*�e������^翖� s�נ�WL�q�q� |J�QI�6m����r�N�.�hA�������p��z��[6�A]ۀ�8�RT�w./r_G.�Tf�k�kt�ko�J]��0_�_��*#��~+��̂��4/��s:�V}�O�ӓҹAn�F����]o�b�U+b[��*7s�&%i��}f�i𝯣����sօ��z8�N��	kJ������� ��!�fL��KP�1cm����=,k��/���9�"�B�V҅�����-���5�}a�:���˟d���m�e�����x<�7�X��Zc�3�ca2����)�('�g�a�Q\%���ߙ�:��?��﨑'#�3ԡ���~�Xp���T�����������`�-�*��q�/6�NT����o�tljOW=Y�o�6�B�ڎjii�$M�wm�
0����R��0��Rv�oY�ڻ �5�n����d��xq쾂ƜN���S$9kjaZhpZ�TX�tC���K�]� L��h�Y?[
[��Qz>�WQ��	�� 1�lxPY��|�
qW���Ӗk�̋�"B�ٯ�4?�u�zu�n��ì��e�F��uY�|AP��C�qw�Q���d��c����K��uۋ�H�|���ާ��j����Z����5I�?��(���b����~�D�kU�-f?�'d-�S������X�y��)�C���Y�{�2��m��ٽ!E�c��>n;���̜n�z�0��0��J�AU�	E�(7I(C�7����sn2�x9⎦&�5���!��3`l{R����%}oa�ԅ�	`Kl�ִ�Dz^�� \�/��P	E��|�Q�����и�A�@�_�vF}��ځ׺�(������­�"y��!�j��ֺ�$�٢v��9{w�
EQ7a-p�U&�_��Z�F�oR�/�+��%Q=|k���?°���-m����*|v��#+�x�� }���y2cf!��QlDPaN���O��P\�������u�ӏ![��ۿ=�oBg����d�2��d��
�r=����X(N�if(Ɯ��P�,{�jC�1:�-.Ǟ�ۿ����S���Vq�'y�IB��������1���
SFY4�9�ߛvv9G ��L#V��VD��"���W`	dV>�G�I�F�H!`��[S�7V"�m<&s����5��W���`M��M���P9�L)Q��=CDwďuL�f��o�t�5[Y������b�/���&��t� �o���+��C?S2��M�σ v��ݠ�.�?��5���E*h�>kE���k�g���6N\��&��C�i��sz��.��A�a�M*׮N�TDC�5�{
R�Q��g�E��28m��5K�T��_�v׻:�Jm.�nd7�<���5�����Nԛ�Z��ZfԌ�~B�9�e4q=����c�E���!���A���^t#�~����������l(q~;4��q�)ԥ�k�tq�~m����TvȤ|�$+���
�����(�=^N&s#����\�j+C��(��ź����92fG������Ĺ�*��}���%��<������Ry�����W����{�sU�!��{d��JrG�(�=l\��姞����:^�
� �����O[ڂ.>�6f'X!��UO��X��D�z��CpHqx$ʢ]PkN�����x����U� �̓���MK�<Ȱ$[�o��NV����>k�Y��>A��I��7O�S�et���׈ֲ�\�swQ�x�V���c����\��,����.g�'Iњ�����"���,HI9~�����8G�Ozd����ЗL��G�U�Ю*�9-v�El�Y!3��� � R��Fdtڄ�{4�t���,Ŗ?���� %%8-himSv��X:�MϸuN���X���D9��6i�%�!JF�L6��(�˄��`�T�{����yG�p�}U�|�_.����B쒊oӐ��	-� Kr�(�
]�B:\b2mJvTǉ����j�S��M7@�!T&!��DK�-		�ohJ�R��7��YȫZ��x8��)z`���U����c��I�#�A{�L5&z��S�����h2��������m���8�(HQ���}joN��'� -="���۠\�piw��%�.�,�����)�O� �گ!f�	��ή�$�E$I��'I،s.}�Gp�؂5�<3Nb'y���h/���������}�~�`�o��@Q`O��G\����\Toc���m2X�r]@�zA�`�� Z׻?�������Nr$@�L�vz��봞��I�@Uc��G��L�5+3���B��lOn. �+��͎������wйk�*��SA�,ʞ��sCB+
�#�b%ī4��NRzO�-d��0<2�(@K;�U�{�&8.e&JY�Q������k���ֈ��R���\��F2*k��U�B+S�E6�\�y$��Lmi�R��r-2�-="K��G
2E,��`߇]n����H"�2�B:�(�&�3�f��r� �4ىf���N�_�i�P%�(v�yJH�C��{���@R��Z����%|�������nOq=�bk.;�H��G�:������Si��7�4`��uy�5�<���=̌�#�E�*���s�^4=���/�m��<=K\߫�q���!�.mi@P�@�f�_�e�[EGvx�.h�֭c�DJ/'���|K�sr�Q�7G�V:��4�ʔ�'�� Y�l$�B)��n]vH�y�� Ӫ�� xҧ�B�\	:�Q]m-C��k�3��n<��:c��+Sh_�j���|�7��W��v!���Żqtz�?����*�&� ���j�>��.���Iwn8>�'�7,�w���W�8��*v+ϯW���������Oq�X�Sz9�>]�D�H:�O��P����<�9�����*i�KY��}�g'�G4`eW
1ޗn��/	�_(�#WT�>8tЄW���0���H7m�����
�ki��7�ԅ��J��Ò�Θu�A�1Rv音�h
�Y@p�ߘ�S�dæ���D�0�+C]e�z�%�Ag�l
'�$X����lU�0�y�ZLda�&�;^�y�s�Z��+#�(��ۖ!r��]q���+F+T'���N!&��o��阞
��삉�=�?����Y��Wd���G���=kS��'�Al��<X��8n�?$����_�Λ!�|�Rx	}S��!����$�Yd�r% �4����'��n �^�9���1��X�D�Cɓ�$��E�I7�!�wX�k�g�,�e�	�(��e7��*�sPEU����@}"Ź�(;
ǉ'&�d�N�(!������4�=y�/��D���N��-T��Z���G�Z���Q�!�Wq�Ջ�z|�Y����`n:E�At��F��v�����i�˪�h���_{��J�
�D�|�4Ųa���=�N�>�1�;��cRR��g�>�#L/�x�E�H	.�'�]Qp����P���"�0w]�%���i���*Еc2#�xc��u�QM�C!�����m��x��K	o���=��P�O<�&���T�=�~K��;���3*� ��O���6T��A
��u���u�ٷ��	����h {��6���{E���.O -��I�<òo!!�V@.+���˒��)��]Ynq�k�0X���.,8@���sMi˨P��&��J/�)�����4&GsT�~�?:�d��N:X{[ה��3f.�9��F�쯀jb�����e�*���
Rf�79v�|?���Q��,����͕Έ�[�46	yӕu�A�D�&g���bx�i#�+�pp�z6G-b�uH�;���э��x��l��IL\i�����M���pQ�5�A��nJuCD` ����<��N{{"��djVm*��	��oi��x�1�j1\��yP�����,��%�e�p��:�1D��iY��S^�"�I����eޏ[A@��_$�^�
�;l��� �_X���d\־�NX���{����^�rCv1��=;�Y���1�~��6�+2�4{G�'����a�3�V
~��ڈ"�k/������[�����ʗ��}��vt�{ao?�J��F�Z�s�o/+JC�������ϵ=!"��k�e�����:r��6�v�Qc�Y�$bc�/k ���p��Y,��o>)���T�������tj��bH�f��ؓ�'%���:���d=����J��WRؽb���qW����
l|1��y%�~�����}������ց���]�	���M�ِZ�9�A�r���âAw���º��d�s��M���4��0�����?��ũaetձ��_���W����j���?��H9���B�b�*�� �,u��j�c*f�G=5z&7���5�A<�9'x��L�2O�N�6����	��䑵���l����- ��\��1��'�Y���dѭ��?t �K�Pza�L�=��W̞�`j�jHg����Z�d��?�-�#Y�Udt�2?�������n(\��u���_��N����x����f����C�)fF��wV����:I�o:v�L�J����Z���S����n��;Uv1@�����h�*���cׄC��i܈�3����Vz��F��]����ap?�§
qx���|�x� %
�����V�KW��>knGV9ʵ1؈g���\���㼐�!!�5w����I����e�i�%�P���80�i�]V�d�4��� ����-�-��3e��'�4��=������Y��n�����0�k.��Z��`�vop�{L�|�3���/	@�x�����:0I��*c�h��6Y(S�&��ᨗ�p{(���+��MS�dD��5���4Q��a˼�ou�pM:]ѹ�&dˡ�ut�r�]��H.Fk��a�{�:,�����"��
�� ��������64sZ����3v� ���UB�j��7WI�3�*.' ]��:�FC$�op��^n-o�r�ku�g'�NW(��eU�m�s�����a�nt� l�h^��������wq���Ӓ�(�x�!⌮3�4�RfKݵ8�ө�W��"^�fÛ���Om`s�h5Bw�C�&8��m���B �ߑJX:�s��Rx3.��D�^��%\��]�E5g'���A
�T�7X���{�e�_�m3z�Y���V]v3H��T솙&�K�_�F�9��խ,+���A0n"N�^�4����Hc�i��
����}�`�aBl��{�m=���q�kո�P��!��~��2���s2�},]�����É��B�"#$���z����\�%�=�,r[JjS��ł���e����a���˿���>�k��RW��>�9G1d?���'�*��a����V�!�6:����g��������P5/��K��ܕ���np�T/����,W\s����]� �n�ZR.����Lh���M=��Ep
q���u{��!X�V�F�3ŝ�YY�����E�ǜ���wjSU��㒉&�x0ɋ$k;��.�+�b���1��$yf��������n��.�0UuL�"����\b����RT�Mߴ�1���/�4��Z'\V*��^.�+��y.+,�,��+�zn�iΌ>CĘlCKz3Ğ���C��%eohAʥ�^�֦<���gG��Y�U�Aܯ��Zl[ W9<�XU?�}�JT�Sf��7��،�w���sl�T;6�+�V�Q˴��1�Z�UK࡛H�0��V����9M��dvF�]JlJwrĞ�t��D����W�Y�U�5M��I���P�G�~9��ɶAd�z����
w~��N��z�h@ FE7���@]c?���W��~b<t�B=6� 7d������S4 ���H��L)�O�Y���@z"B$���諸�|sU��7IB`_�'lu�ޭ�R��8�`k�������F�7*oOS���^R��ɳt?G$;:�^��Wތ���V�ý�K��с�n����r��5c~x_���>������B�	��dԫ�N��,_����"L���
�%�k8��+)ڷ�[o�f�vLަ>X��x��m�8����2�&�QzfW#�ـݼ���i+����j������@�8{�%��R��#�w@lN����(���,kl���)@Qp,.�C��\Yy�^m�kj<'�D��#��Y*�"�� ���ς��C�<i�d�$w���5�Pn�7��`<]����GF�A�L
Ү��s�'��*��3�����r����m0����&{w��{����J�>��Afv ����u�T�Ki'*B�NS��X���|�mˏ�-��d>��40�7j�j�%���q���!�I��]T�� �F��]Q�g ����92g |�
�dq9}
ťB�.Az�U�'*�MO�=���F9�2$6�o��d�&QA0��C��]��{J�����]Z`���e�6�4�cʈD�w8>�ٯ͔w\���H����)
�$t�E�Y�]��ѽ�jK�kD��}��T����Ӧ"B���70/*��1t�F_
�[x:��n�n�t�,{"��Ŵn�9)r��RR[k�����6��[
�6� ]����k�M	���<J&���L`xtқ����
�����,4@����B��T��������r������/�8����&����-�I���cj�[�><4|n��oϣ£<���Y��D,薀ړXH:��R�۴)U)Ι����m�ܿ��חM�N<s�yqXb���wr���R��6�����_v>� �еK��!+�_��v��ө�ْx�i����̄���rTZ��jD��2�Q"��j��*t�F��ՕE|;I�#s�&&M	P��g���� �4ښ9�5p��@���K�D���w�WSO�|�`��D��m2�îa Z��=��E�Ks6��f!�gW����U;���R�X%��F��wW2�f:��%MbV721��e;�VD�ϙ�@����2Va����Zd�t8`�$�|\������>�h1���\Q���ȅ{7�$�ڎz�8OH�E̤�㭯m2/lèn�n�+n-�����1:�
	o��B��I�V磒D؇�t�a���(^ƼT�ͫy�h��s^��آ��q�����lӬ�XM�G0H`b�Y�9̙{>Xj�_5$��T�?K��[�+���%PԂ�`J���k����G�޿$v�6�,W�넭Oٳt;��B6:F����p]�e�z���ZY�Tz?5��qM����~Q�s�A�8�H ��D]���l�R�P!��cV�f~f8*��E�SP�0����R��Q4��ЎC}�T�?z;����sX�a��ڷ2�qϪUZ�BS	�֝`#KE30y1�f�(`���?s"�y��#i�z^�0Cs�2����o�6�F�y�vh����a��(1"���h�KK�.ݛ����G��O�~�j��I��>�E�E�E�p_O����9 v���g�ܗi�o�;]����Tw'{$5DB��.<w�~%歼2�Q?Ȱ��bxk��ͪ��V�gQ9�nm��fL2�)Re�������e��h ��`S�X`�vѲ]Z�κ5���vvJ���Ĩ{ܔ�w�P�"L�����5c4#�� 4��LJ��o ¸e�T����G��f��ÿ����=�����d�W�/�����n�x�]��w��MM�IS`�����.����T译���1n���#{����H���\y�g�Ϩ��H_��R���8U��k��C���,JRq�	Ҽ�$*�6trZ��7joQʆ�w�{��?˷$��O�ƨ����[rS6gg�tu
*�.���C�NpL��9�c��NG�Z�v��ZN�g�JN�z[r��4TrrOm�P{�6�n����ooC�y��U�C� v] ��[!zF���4���w��<<��{�qB�Xu��zԋ��8��u$�	��v^�;�I~Z'�v�|��潮��;����fܝ�A=�'�噺l���tb�$ �� �,x.��2y2%J盈�J�Q>b��L��Ѿ�,������ˍ���r?v*]�ו&�
�<�ѿ��k@X!����)�6�lf��]/�FKh���:l_�什�^�
����'=�c3�}Tq7/�p��a���C�@^2��J˗��|�Lt;��6��1i�v!�`$o!����4���0���ێ��z����!�\h:���L�I��'o�xYY��9��,]�p�+�fP$��)C��Lé
>����3!Q�%�:���}2�����#��	��$ �7`x#�C*� ����Ơ~�2���]/%@��f��ǭ��y�;�GmVg���g&i�[��V��=M]s��R�6r*�w���ٻq��k���C9G��/.�9ÄFd=~0T�	���C�������b��w+Aސ�M���+�*݀)��a,?�3��.!������j��@�b=���&�� 	�N��2���X��Sی���po��Č�3�LBKh�������{^5�� ��?��V�?�0�E�]I�Q�Q=ڏ��P^�����O��_�s�]*��]ˑ4����^��F�	������m��,��B3Շ�~$�}T�<�G&��߹��@Mυ�_f�B�en�0bB�$���<� ����ZH8�����������}`繵�0���hy,e\o�G��g�/�=�Q�}WT�k&G���w��c����<���;/w��(�5�U݂�^��X����v�N���D�o��1ो��א���v�"h�R# "ˋ���z��ނC����"6L����]��i�)uq?�`���j�d��3љp�Ƚ�����=�۱'L+�2u�AJ_��]�����M�=���#�a�yF[N��D{R��/��#��CA7��&�8�rz���V��|�V�N�)�b�?u��j�CW�rBl��'���	�\�j�Li�R�T�ɮ8�-p�Z��t���*�)�e�WA�h�S��� �_����OVS�@W�±M��Q	�Nyܨ�?2s��Z������?Ŏd%V� 2i\䋨����-&EG�GTn���qa	��0Z�4���N�uG�Q��
�
\`w�m��y���d,���g�A֚���/�墆`YsK~�k,�H���0)���%H��K&&MƔW�,�N��s�=�5L6�7�[eOU�c��n�$D�!OEc��E�,Q���#��o���"uPe&d�V��E��	 ��D�������vx=���硆���a��h�H�>E��ǅ+�>Ђ��J�CH)qA���y��)i��|�GݢBC�p#g�\H��g.�	��	D��G�����o@��3��jӟY�P�ye�C�6y\ �$x�)�F������Y����c�])f��;�v*� �rǨ��-��2��� ����}��6lb�n�E�l�i�=���e�&pu�G�;�Ha�B�S�<X�Y���n-�c1��a���g��i8�!��[�s�A0���qr�z]D���6��6���v������e�Qݼ����n��̀�Йȵ5�>[n����,2!��D������b�|�]�6P�o�,5!Z��m�kL��-��^Y�ݒ�����6�s��ҧD����;Oq�����_�lm��};�#әV�mZ��#�g)�a��@��r�	�e�����X}6w�"�
|22����%FZ��(��5�m�����k���FP�ƪ`�3�įq��~Zo�/S~��jO	��Q��T��O�];�c��2PAfZZ�a*�y�\�u�[�� ���
u�U7�@��l��_Q�Z"��@C���O;�t�2I��Q�d
I��w�@�Fl׈���ƙ(����_d� ݙoN�j���d|����6���|I~�3,!��UV�oi��q끺�{O��'�EA��`��h]ը%�Ho�M�t��A),
D�ˠ�}�TޕUD�?3q�f�9���A	r���x] ����7��c�g�D[x9�/JX�3�S�W��Ԩ � Lr��?��ǿU�1����V�Q��o��$�?�?��3�GB���������3�J���(��za�k/h��$��_}�n�Ez3ƿ�:CKDA7椉��T͟3h�Kr��㻾u ���j(^1�L������H���%���(�XW���gd�v��Q�/��7��D��b�w�K�6��?e\�,�6��E������� o��NCj�A�^Oݠ([9<I?"���EK����,��L�=�a�q[#��h��ް�߷$��H�X�Z���=[���(_C��	�5&�u�u[g�݅������@�&�ӭƶ>���y��IG�[`:�E eQ3���V�ˏXw��E���I�����b�
���P9o&��;���X#Xܺ]g�}*�Kʵ�&^:����9x����d(j�̨�Y�M��9�i�����K�2�²`d�r��VP�_do�vf�|�ܩ�%❽�	�3��B����;����@�9��G���nɞ�x�Gw��hե��cG�C\�2{o� �#�#^�.�ϱ�ܳښ�{�W8�b.�i��1����g���K}�N�%�M&NH�~�K$�NwhL���t��~�+0;P�5`!K�ZE�")�с�d���cy�E�|G�����ݿȦlS<^�|@�eJkG��'3�$��ç�%�*�	�l*Ϙ�n�5�.���9}�Il�-t��|�ݹ�A��s��'�8L"�Q2��m\]D�Y�_�����^�E��#=��'h*���^y�z�o�k�a�_�c�c6�#�S�I�
>�N��hd�9�T��g�0��^=�e� �^��m���q�E�0_\�;T�����)��z�w�*��� ��-�ة�c��.IW��M2���/�q>:�b���l�
K*S�ӥ)����7�O�՜HJ�j�S�0��Dd4i�{aI�k��Ʊ�C�������kdKbl�ٞ���s[���5����p铳�@O���Yon���}1��(,��!�Ͷ��/��\.2���� f��.������K^)^�\V��؇^�~c�>����W�k}��A�f��D��Uˤ���ڻf:b��O���R��-�^S�ɿ�}��uE�o��M;MM���N�I�M��PK��m��:r�og���\��w���8E��(�i¸��芆��F�����vо*m<y�v�D��	T�s��������HY�57p醞C�Wk��@�������B���� �4Z!_���n����	1L��:7c�|ܬ�:Ć����H�٭�%��TvQ��z#<P�����Ӛ�d���+����NR�Y�h���S�W�j :V��� a )���z�*�8l�m�h�f3=|F�O6�t�u�:Z~m�x����n18R2��<)tHc1��F�x��^W�����T"�>U`����`N�
)���� �u{vF�O�����d[��8-��Q�w�<M�u> D@�~w�}jң�)�3�K
w���A*�ݧ���KJ�J�,�;�o���'7�V=ڵ0�v9lM99��io��R��ҟ�_gX~��ǎ�9�&�OY/7�:�H�NX;V�Q�K��&׷b�W�x���:#��׽��L��2��6=aP�li���y����@�7���u�����,��j�y/6?A�`���P%�����P��"��,�e%�g��
��9^�k��a���̹��6E-�dy�*y�;o�3�D7��f��3a��?�}�`XhR�+�F�9��L(��X�\�AI�2,ԖԦE;�t$���S�?*o��gC�#�q��&��!�����E�J}7t��N�o�y�TZ�4��&Ӭ]m<r�E{�a�X�xv�޺��q�I��>�0Wü�:��F�%!�������i��|Ǐ[Li�&��H�b�͔�A�M����OݪJ�k��ѕ��
G����L8�Y���X��s��JU�|]�3�r �O3� �� )c��!��WOiM���g�kk��jn	~YgR���{zI����]܇���s�3��E6�"�譈���A���W�:����F��
���d�R�7{�����7�˘�K�ht�a6ڒ<�uM�����b��c�6zV"{7�&�8�\)��%�R�jr�ܺm>�>$V���wS�I[ʖ�锅�f:.S٣�-�x�T'��d�i��UǀA�G2�\Kb��H]�9��a�n@E]�چò䲻W	��!p���K�^5�����?��뛤.P�@"<��J�ٜ�ݵ��4��	'B