��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%�׆�o���L�^���l�'�7U Fi���-�ae�����$�  Q�Z(���Z�ǅ��YX�Յ�n����M�r�%~&O�suQ]y�m��j�E�z�TB�6�-F��r.b�{l�O5��C.�n �a�	jy2��<��w�o_�k���,��O����u_)��i�j/1}�:ZzIJW��I<^���X��uIO���BRu�p4�K;�uӗ�T:�����fiZ��kנ�G�ǑiP"��z<�,���^�,�_�%���4cl��F`6�]��ʆ�-D#-�a�jͿ�����v[�)'i����p㺻ʪ|p��Ɲ�fD�#�C���j���k�ې�Y& hd�v���8�`X��>:}����`p�|sg0a�pq�K
��eW�l���j@���E����V�?�g�T�j4x�*I�����1��wL��_�A�遇*��;�e��)�_y���X'5p�����"7Y(h 0��L��4[]e;h;,����w3	jKfw{��F�꩹���s]���Z�`�A#ᄖT�Յ(͗"���ԂR����:.�d�ysG�p�9��ds��_l4ziK��N�]��Jf�s.��Q!���[���L�����J�)U�r��E2�&�
�T�tQx��t"�u@)k�����f��sԗn�X�j~n�z�^�H��-�'��k w�J0j*�j�c���?�0�~2Z��]/�]6 ۞���U�:0sj��&F֧��3�c�Y�>�$U<c��*)��vG���u�W�2Ǥ{�Z藻�#h�K^��4���q�Q�	�f�-ǝc�}-�j%U%TT��`�yI��R�˻�Ǡ��_O�$�������^2�>���r�z������y�Y�`�w��"t¶1�mVk[ �<cs
پE�ͭZzǉ�0��5T�1Hv(�#?:�H�]@��Io��3�U\E��B���_�q�N�7�Q�[�B����2^�H�'��󺅎��!R�d�;���G� ��,�?�,�,ӑ���=Jf/'^��%�~ˍ_��w���K�"wE,(P�����uͼ����;�jK�Z��;���A��/�d0j��M%8G���{��2b�C5�[P`�v����8�WF�b}I���������9K��7=�-F[�x�oX,�hԏ��%�~���bc0���	���#{�@͘��R7�P�I�p_2us�4^�\v��ޅJ�m1���5O[��s��|BV�?���b�3���
�~��G�dPŶ��n����Z�g�?�0s%�`l�][����UJ(���-��i�qm0�t�ւq�d"KK�_�]�'�!X��x��X��_� ,@a���'Ā��;��H��r�{�������T��OO X�s�v��6�9[���RA�[�@�n�}O�J��J헮'��#�U�%lLL�n�l��˫��M��x��*��P�2Q���vm%�mYuI~D��(����q��]Ϫ#�F�bs�j*���#�%>��j��8J�%tt�NX��k�8�9Ԕ?w��qR�gGJ'
��TC?�h�x)���r"�kFBן����o����H6 ��N���ĭ�����\�c�F�:�ٱ/�Ha�譠��+K"θ#?��"�Pk�?������t[��Q9���e �+O���T�������4������i�B=��}�7��*fJ�xyW����?����Z�2�D�j����u��4�3-{T�S�� !�=͢�Ey2:�s�֘�W㽻��/d�e��6dx�}v�2�	*)N1.˕+OIh��)�S�0���b'\\�c�ϴ���.���]��L��"\P~B� ���f�q��<9�?���"X�0�ڍ3��qsV�;��Vq8m<r�q�F��H� [��X1�.Y�6^���z@j��#K��3	�,�a���7њ���+#��'���QR�c��*Mج��k�SS��s����D�?����%v�}G�3��]Hf�5$���Ѓ���u����A7K�RJ��ȓ=�����bq\:������#KyxPkԄz�q���i��4 �lR6W���-K��+|�?}�W������K:�'��T��.p�6#3ߔ9S?��St���Z��0�Z
�G��)i~?Pq+?R�*��2�f���b����[���;��=4�ucÌ�ZX��h@A,�YY�}0����H M�����	[ӊ��A�s�l��dyR���<(&���P����������́���CL���N&q��P���E,*d��vw���6YfxW��~����� ���/M?5��+�eML�V9����]��E�/����IH�.����[0�E.���+�'�n!���S}���+�m�1�0�Tk]okϴ�t@P��|z��7F���x�xY��U?"s�R��C��=?8��{ ����bU���$"��8M#P$��}`�;�7�?�\�T���$h�0�>�]��2�Y�A���`8E�x��n��]�Qxzь������fU	��N��CI�w�X�g`�$�b��a��	:��1cK��<U��<⼩��S��Mڌ�g�̬�9]�*�5Zݡ�5ⅾÛQ5�n2��11�4�]<���ȌBU)ċ:���F��������%Ѡ	bi!u6�x��O�@��*�v�r�թe\T���KJ�Q��@�isը'tzz���0�vhЏw�?��p�L2��
��"�┬2�RF��`�Z���u�3� ��aн�&����UB�Z�^��!Ͼ��"�G�y��Hգ�H��f�]f�����]��
��:��p��Ӧ�+m���.>*�{�&�H�jM�>�¹l=(S��2�z�A���OD5�=��qkI;���L?�`�]�B��~,�%����1�9{?Z��R��kzƀ�f�#A����-5�8p�l��,����
~3e8h�ı��x�H��#�-Gq��|I�G������IH�#%Pe)�rI��v��sϒY�e:,�����O�	1��I�o@L�?}w��=x9/m��Ǔ�~��&f�^���}P��o�ڐ� �U���r/��i���-^#��<�c�_�X&�0K��	���Y���
�[5�5�f���yk��`*�%J�+����M��ʪb������jI�џŶ�	�'��
�f���㯓��_��TFv��W�_Z�>�4�jd��C���5W��.�F;�ƭ�]EM���O�n^YG����Y�EF�'��'��6[}tT�iK�}�@�d�7zk����r�)�����/�!�
�5x�����4�E(��R�(v���Ưj�gOl�Ŭ@�(�]8�T+�񵛆���u,�bGȄs���@�������[ ��i	u�|�F�S4 �jIm��=y����Gս}�I�>���i����!��hR����%�@���p9h��4� �OU��b��&�i��A~��P����^���
�?��)׻:�Lx�,h�X�"$$�'�Q��Ÿ^�e��<��Q��a�l��kPn?�w.�q�Kp�.	8a�Ȉ1�˪��}]�!H_A�nS5��/i��D��c�"�~-���i���-�7�e�b62TR���Y�S9?�GZ@/�ř�D���}�
֋����_-��V�K<E++G��<�p��?|�����y���/�v*ގz�tB���"T�c%��Ba{�����m)N`,~<�Z�ӛ�%ChIH�U�8=��#���v-��^����?�7�a��	ঃ 2l�^��F��@��~+6D�R!d��W����mR:������,->��B��0���e��d&0|N�*�O�?Q+��5R�F��n�G�\!��ǳ^����������V��֠A�Y���D�z�N��+_.2�v)���'��i�3���HN��a�>�.�5��Pw�rdL���#�w)Q��S�����c�GE+����ޱс��w�n1�����1�z�ÕXBR\��{��7�c���;�N�9�aM��q��y�Я�&V�b	���0�qy `j �@?�\H��Ki^��_�K�l�)��b'���o��V|V����1L-� ��˺�n<��}�'���I�%a��ڪ.
��YOAоR�����îH�i�:�rt�s�R�R9E�����Q��4�����@Pl��H(wt��<�\�}��~�\�]V,�]���]��ޙA�=2���ׇ4G%L7�w��ߨ��N��b�zNd4]�3�*�Eu�,��{��u��2t��m��T����M��"S�?0��B��Qp^%=3�u���딦�O1o,�c�� c����f���/�"���� �aey���m	��ƺѠ��W��;ƒ7@lZ�����;��=��&���-�8�*�;��#�)��< yB�w���MT!��#Sg�@I�*+���g#�����`����se���<�9+��Q�������I|��"O�S�'C�h���E�	��)t���1��ڠ��p-[
^��ĚTx�a��pu"�3�����t�x~��H��P�Ty�^ǥ~̼�aB2S4$��:��:���g�����tM~F�h�>��G޿�߄ÆϪ�	aB�2z�:L�w�e7~�y����g�-�8��- �?6�&�2`
�ssLpRv9�9%��>*ގ�L���<\N��IWiG�d>~6�cQ~a۾5����x�ikYQ�쌽���I�-c[�/g���xK��IN�q'g�fe��34l���~�<�=2GW*��6J�2֮^�I��S�"ym�7-G6޳��A�A�!�����JYϱ!������g-���C̉�tK��S������%�T��'$QX6�C�[�4�,��T��v{��jU-��?у6�1��>�]6��S�4���"���	1�}�����A�e
"���	�B�'�V���1��_�9�.4��S�k�D�f2ћE�
v�%#b:܊����C;� R� �LwyP������$�.��e���%�?��#��Z�f ��9���O�=��6I�L�02~�_�c��U��t�f��]w[��.��*��H�G*�w{Q���<�����A�ۼ
|%:�č� �ħ����{��X��OQҾ��j��*�Yng�f���K!�(2��ܤ���\�+�Yک�f�j>|���Hf<����U����bD��o��зZY�F*���TI�<�#y����ݿ2A^y�6A{ Tt #-�51��sc����}���T>B4l9��ݎ{�38>"�M��2׺���lJ%'�l��c�W�ɉMu���a�F%8��[��X�<n'���Pz4��:���d��G4$a�C%H5|�F������ ]���H�qr��j::�F¨�δ@m�t,���g �;X �O���%v���hw�uF?����#��zZ4�I���CY�t�q��v�"H��-��f �Ntq+P���68ĕ��7!�D�se��΃�K5���*y@�!�Y%����:2]�f?�g��u����^�\Ι�4�T2Gc�}�/��P�>�"�H��$1T�ҙ`Cl1@�jEl{��^����]~���-^1�&�:��
K�H�iۼ,��rw�Aa���$����ҝ�4a_�z,*���e��1��������( M{H\)�'4�?��H�+�O8[�W ���&�������X��һ	�s,���N��G�Pn*��p�fy�r�����Qg��qwϦ����0�}���&7Dԣt��H�����qE>?�(�K�y~�cF�`��S�W�d�:�[�Z�5g�JZ��д���/>�W?�W�9��:�/u?)�,P�&}�K�Dk��"}.�y�8o�)��R�'<�t�T5L�X~���K0ҝ4�-I���+�@�v؄P�F����1=�q�BT��Sq�N˯t�ʞ���W�:��0�B���pv��y:���2��π��p!ٱ$���W��u�r)֢1�M�U�ӥ�X���xmG|���i�h+N�!�L|���6� ����Gy�%���10�Iȅbk�?6;��zvI�'�j�i�X��m���F���}���"�tf,�T�=���	��u�z~0f˷���9]ժ,$J��[C2��<LkP)�P1d�r1� �Ē+����.����`���#��<��NmNЛ[��(;��[�>&1���ѧ��>���^ ���pw���Pc���5r؝6�A�RW�}u�yY��o�`�/'	W��u�?�;��G-5s�&����U}!D��ZfJ%��j�G���{I�C���x5	�bh��[kjO1z�nRJ�E��#��c1@��I��5�%�p|�;�U�V�mIA��<`�
�&҇�0�l�d�|1;���	ѧqWX�^-P�X[T;�SOPWx �G�k��D�f�V)��2�c�˟�,�ψ^[.|�Չ?�����2����H��9t��u��~���7�u�IMI7�ܹ�l'�w���v�"Q}HN���"�Y��[W�����P���b_�(y"Ǿ]U*�B���x��|�8�DN�%3��W w�
����
�|������DT�2��0/�i�k��!�8���V��X�9߫)�
�1�c���1k���y��{�,�
�0p}���Z��ؕ#+���*����c��XHw��s���\#3��'l|���ւ"�UnB�Φ:k���vk���k^��9<͵��No��.���oUE��	�X�cF�	Al+r����|S�L~4�H9pA��<���9�GE���}�4��q��|��uA=F�9}�9��"?�@&��d�G�#�_Ň���k3�e���KN:���D��2:,��"R�Քr��G@/���b�G@�AѪ.?QY�OGH��=4^�!�Mf�l1��׷���4�#��]�`������}l���z�$fN�;�QЭz�BͨdP�����c���ЂP/'�]"Ps,�a��b$�Zݩ9�T�9^�^�<��LZWI߳�&ߏ�:"�x��1c������H?��~����O=��2�SVv�C=Lk.��H�j���0�9�SG��^�a�p�j�?/3)��#Wn�d�..~v��<��5��g5��?������+��B<���P����7m�K#��G��?_ʓ<�2]��Q!C��fZ#��K��U�L�]
�u��|�PLO�-=�W����nuՒ�l��a�(d))�$���O{�;�9oY�|\�%i�V�~��^���L�^�W�:Z���x{��mC�5�?�KE�H�0FS����?b��o��7^R����P��n�&-�����e��������k9(tJu�L���90�6 R��i��0���ȪT�6&gmiD�_��8×I=RH���1���,e*i���~�� A$�TO������ �5i?J���F��	�6��k0�H�?}c�?M8�&&[s)-���0̺HI|xd/�[T�u0��&�S�;v�z���/����ؗ�ҿȂ������эпP�D��-�}��ꘖ����t�P���Zu���p��?� �3q��[sy�L�h����O���7�%g���u�Ҕ�F۳�V�j��]<� �Lo'+!��vc�	�p�2���_*�@�H�`�ɦ_�0��7�=�_�K� ���܋�4����W�r����א��*e�w��7��(x���=����!V>�	�_��+s�sy�d���X�FD���:�5a���:Z�H,e��[4�x)�m�t�)E��˃�<�1~?�޸ޟ�*�<���i�U=��\`��9�mh6���n��h���k��M���  8��罽X�`NbL32^����-@H*]K�
L�0�$w�Z�NLN����Ea0��g�d�	�֑��c��!�m����/���VJR�)��l��O�m/�9� ��c$@�#5���D����y��&ō�,�&���X7%��G�5F���M<U��M��qW��������=��/���$���='�$ j�j^�_2�k��^�|A�C�ml���ާר�x�JK��7�q�6���l|��c��祶����oe?�0G3�V@M�x���K���d�e�0I���DJ3x�4\��ث�d�L-\��}���0ݤk����!�[�65�<r��w�W�G�(b� �֟���N�_�����>�_����(�rͶ����@g]��������W(����͛B�+������<K��@p�q�'�Q�?Y��9
'��ƂZ9s!��X�0q�kZrYt��Sȉ$��!�4tH���9d�%�s�045ɱ����&��o����$%m� �J�����$j�v�cQ�+���A}�3�� ��ܺ�PJ��F���Q=�u�b(��;��5�o	�b�]wVQ��๵�� �U^�A��y�7������a���E����l(�c�@^�`��-WO�_��ɣ�,��$4�V�<����ŀ&~HB���4T=�b�{A�PC��y�{�U��[U���v4��O�m�qӷ�m���w{�F<.l����3j���M��;X�VJCߗض�ˎ��$�K����+�$��Ew#{��ln{���<"�˘�8z�-�n�G�5>�S��F�d%��)������Z���(�`_8{Tw���l��45�f���F���7�;g����	�u����|�s�b��>���H2�c4���H1�猝�m�γ��Q;DJ���#V`O�i#U2HQ[F��ł@���f�MK�W�?2�N~-��J~(��,|�MN-�3pk MYgn�m�Iu�7��:@o��A'��*��@�2�*O6��c���ʙc�C�� ��Ț~�Y��Z��"T���#f�b���"�$0a_���t��p�Ə��CJ}�������XQ�m���8���`׿��C��[3�n@� V���DiѦ�[��Y�� �3cW�F@�W����+4��q�5� i���&7�P�Ϭc�{�u+����C�Z9��Qt�]Xޑ�>�̅��$0r����T��=�d�;�M����ɔI�#N`�tS�C����m��P��n%S1.��*���z�A���`hs�v��!���b� ��!��.?f��|���K�'s`�:�Z�t=MU�G����-�S�?-��}�����Z ���_����0*Cr��J����떨18��m�u���o/�I=�����MA�"�� z��c�uEc�/��h�����Ut���Ȉn7�������5ľ���1]
,�����T��_rٍ� g��B�my��.B����ê����� �{�O��-O�Kg��G48�߯TOL$]�N�����`N!g�o?��'QY#7�6��6�E<��|e�! ?��A'�SI�S��T�5))Z�7PS�+Fυw5�*�N�S'�kyZ�!��oP�*�kn���oAΤr�������v�[����/8L�F��������u0u�N:]% �\|]�����"KGK��X��1�b=$e-�R�У�̈́�;�vo>^���PJo#�$��ba���6�<�[�Q��S��J	֋޺>���+��ገÈ!BV�A(N0e|"aE�C�t8@=��BaطIO�F"yX�l@��(M�[���Jɶ�Ihא�� ��<�]L�I2�N�MH�kl��h����}2)�	��Y3zF�����&�P{��/�R�r�l7��cR�*�Q�ղ��]�9�vg��C)m����F�x�P�����;��v��"+S�; Ǉ��Eu�M)��~z�������ռf9,5E������5\���G3h'&���y�br֮[�ȳS�����ÿ�fg{r�#�!ʭ6q�
���]���X�Py�_�0�+erm��b| ���gv�cux�+��K%�93���	2���{���#f�f��}O�S�CQ�JI��BK��p�R��r����pX	�'���T�$
�$�@Xe�F�s';ts�DF������:�R��AΞet��T#a���<�:�1���(�MJİ��M�9��ODn.�gD�Y���i��8>�S��vF�5M�~�H,W��L�W%�ި�s�o�3�-�&����|h	�F>����cve����(�ʧM�����w���ލ �1-�� �S)���?ܔ8�(y��RN����¸��0�R�Ρ�<��8���c�L3�����E|�nZ���)N�΅��G��{��t�Z������zn�
9K��D�q�E�,D5�6̶��٫m�g��*���k�y�/�O���N�S�G�˯�<g�9�� !M��E3���5�EnZ���V��GS�6�CtB�D:��*��v�X5*\�A1�=L��';E]/���YJ�Y�]?BГ֞���c�`���/qK���{|��6Q�\��R�+"��<�^xˢd���Yٟ��dE�A���8�+X��a��������9�R������M���:%�N�݇��oBfQ��`�߯o��Unl��P�GMh��DpE�+͏KԔ��3�vM� qp��N�گ2��a(��(�A�^P9Qq��L�����r��0���E�ޏk���Nx͕�E���S�Z��u��]Z��Hn���{ ��NR �&-g)�&�T)Ӣ\#:�4ʁL[z�V{F�̞�����i;���ppi�����KS�x���2,F�yk4m���xf^�YH��e>?��������]��V�j��*|�k1xدz�A�$?���ŊS��q��p�2�J�j|e��Nk�L��@����~L��
������PaΌ�zL��0�oq��C�bç��	��5}����-�:tC+�&�ue����#Ыm�z�\��C(g�!���,�P��ӌQ�T���KExc����p^�(�b��w������3Ԏ������ĕgS߭�!Ŗ�7qD�e�uLfAr���
3�����u�|�b��A�؁R tK$쯩V;K;��v�ʹ��������?x�&�g���O�)�f�$�"2KbF�x��O�dusx��3�,���OԩN�씂 ������&����	l��MLQ�b4>��ֵ�5M!��\�t�ۢYi�#(=b��n�9c�#-�c�<f~Di�������9��}ԑ����@,�!�;%j�i$¨�蟴3���cL�ߡ����K�;���<r�O�S�%�M���Rbd�Nl��(f�������:T�<���>~k���H�ُ7��%�T�U/t̡j{�Z>O��6���A��骐�U�Yy�eP�'��3ĝ��ґ�4���B�;ߍ�+�Jh)k�
��׆5Rm.��;Z�#����	V�ؤ��_����^w�rb����D]}=}@ǚ��TZ��S��;�M.��L9�o�YoV_!��|����2�E�o��ʫ���>�H>�o����> �1@��G3��,���ϵ��"s�6�>/� �u�U��/أ6�鐴�X������|Fi�'�X�h�����?d��y ��V�hD��f8?�#��$���.�/�Eg�b�q�N�.�_��t�X:~Χ8�*�;����4�W��P�o�����32o�[��D�����z�y�"{��U�U��@�5�o�)j*��x���rQ�;e�)�}�����:�H�>�LG
�QN󿌯�P�1ǟEx��i��Aʌ��{;�"cU=����NN�M���<��		��Z:��� a����?q�=o�i�#�Z�T ��*�
 �O�2O!�
�SF��c��e`�K�z����Y��m�8������!W��妶�W5H�-��E݌ĝ��av��eM�	ǜ�X��0��v�\q�Re�ԗ*��k.o���>?:ck��]o��[���\ �o��A�w��8��3��ءQ���Ϊ��J<��7��V��%�3�` ��1V�}�� i��8�s�7�Q����QP�Z�S��9�z������@��`x�I_���r��<1B��r�~,�dG	��פu��2v�F@?T���� �:�Cr���I�yC��O���ђ���Ȯ߀)Pf�EA���f���͘��v�ѝ�M+S����__�֙A�Z�%l��3�?��nkC�0l��� 7�a~�g��a.�x���1.N�"XqC�	>�5���I��*cme?����QQ�^2�7�^x��w�-���	��Cai�)��y^k#jbۧ�t�A5q=�lJ�;۾�M��Ʒ)���_[N�x]0w�t����,�Y#�.�4[��HU���ߌ��*̙����o�2����D�r��|�z\���9ObI���0��B��xBp�D(�x=���&��ń%S&�	܍��[ê�]Ԯ�DE��\�8*��i­8͔�Pl���W�.{�6z�vno��-�H�1\�HI��+s^k14`坆K��O�ā�.&\�97��Bw���m��Q`���y�^��ف�����B%��7"���Ҁ�l^�IOq�F�h�$	����,�T���$���������fɍ��%�%���}5�>#,Ȗ�O^��Un��h	݉6*�Z�]��E�T�|���KA�L�(�칰|�^J�u&����mm,� T��/�0o�����9|#K ]#n���+Mb5^N߅����-3d<���=t�K����f��/o���u�Z0}E$zҰ�����^>��1A�,A	u��\I�r�E�#����~�0��������X[��ʠ�؛���# z���w`�Sy�)��+F���
� ��A*�bVɉ�����s_\���g^����T�Ճh��r^.Y�S0��n�I�|�P��7�l��}�ܷ�;���(";��*H&��g#������-���G��)�/���V	4�h��#�ad����=�o���P���X4E�Oo$ρߊ��B��՞:�tŪQv��Z�����|W$㬗��>��-DM�~Z�7i<���j�ÎN�?i����j����R�ˢs��= ��wk���;�[��	*H�'���#M��E���q�>N}��H[]/h�X����a͇��A�ط�x+������ ��B��4-6�P"W,'
�2��Y�TZJؒ!���o�#��XF�>�oȹ��y	o��YY�k�-����7N�x5O�Wʸ��R�,���D�k������y"n.��9�k��4� ��˓%�Y��������1\�n�o����M8;HJtΊv��������P�}}U�W�����)kF�"���K�E�ͷ:?Up��t�6ހ��gjŵ�Z��2�}������bu��$F���^L�(o|��wʽ�B�.~�ؠs�c4u�`]����?\W��,�H-��o�̄�<��\�P߁p[Ku��]�c�����(U�a�:�}�����-'<S�W*�&i��鎙I�i�7�@u3�p������.�ޤ�٤v�3����aR&clU���{l�:�:�g{ox�&Oخe��s�;���s 4�@�W��T��`<�c90�Z���/�E��F�I�bY�X� U��y�RK����p@�	X�S����'�����==�ӑW�<�q~�fkn��ی�b�]1�)���x`t-�����|�U�-��Ҝ�$r�r��׆SQbSQ��m�|��?���ǤG<�˷ʒ;f�G_�!�����L�����͸a�hx
��1���/l��D�l�A�c2V����B9���>�*c�I��x����%����Y��� �v�&� 7�K��!|����=u�w�'~��ЅT�5}"������'�N4�8�<n2S�:e�	0�
i
�u]d��']U4��y����Ռ"�;�&Ҹ����i1i���jP������Uϋ��Ϥ�)̔t��l���l/���ogP�Z˭�򉯦U��W��w�\�!��]�( �����߇���~fV���R}c$;p�ԃ:)���tK9�1I���5�B�U[��uM��1"A�r'S������0 ����-��d����o�|%��r*�1���٥�9��=d�������$G[� t|�K��{ C�pD�j�Op�	4�Û
L-�"� +�Ih�b��4����`/��R��p��w��5�2(��OsC�gcf���m��_�L�.����5��U�N�x��)����~��qp:�����9�Nlt����2�8�gU�;.��<�>t�oF����Z;�]�$��3� �5lx8�����s$1���
�E$�$��}�х���)yB@�o$r�}Y���ི$�l�M�ەvh
X�<���`\'C��'��|�{�T�26�7��;^H�7�o��B��[-#����<Q���ep����
r�-�ۨ�����4�I'2�/����-��� ��O�碪�Q�q��V���X��5w�є�^�t9m�d�V�볧=rh�բCO�q���$��5��F�U��a f�h��)����w�YY�┵�(ϚJ��]F�}�I s��񝱼]�!F�3A8�/��SV�v��M�&�ne����7��F�1m��M��U	�T $�;>���q�0Te[��`1�P���s	+t�J
wT��I�~��+r�:�'����E<�>��v�:�%����G��^W�@���_BW{�ܼ���i���뀙&�d ��7�2	%�Ťv��x4�-��	�]�����A3U�*�Ԋ���hp}�����)�kv>D��}K��eTb�k��-�#]�lT�����C�+�/i�	1�̂+��"�o�,�a}��h�����~PI���Mp�����ٶ�y��`s�}\�y��:LCR���i�W��c��=�9�M���]¥�d1�V�V�o��\a�
8N�`;�]�e� �tĈ?o$^I�mS�	77qYY����X�8�!�z��0���/�h���"��[�Q"	��7��)��fI�����Q)^/�A�q�W%!z��3�������@29/����T�[u�K������c�n}gYV9w�:��A:�5]�~�aC
tj����n�����<��R�!['��o��K�g�t��\�c{[�τπ��iY��ϐ�Q OR���G=^J>X^ju�A;R��F�0��wf� �G�yw�<�A.��H��0��#�/V`+�z�RS��h����y���v���/��8�h.%m�8�Z���b��'�i!�0��
�(n���
�TǴ�d�꾝��	�gv�r���.�1A i�&OH���%vrV�Yo0�Dc�3#���:�=�� ?lÀ,*i���Q3@.���P�٤ʶE��Z��N8D��	Jk�.�ٶ�[�d�KT�J�Y��⡗�>�7��Ń�����I�G���>�j�s��W~h^�������۱c��1TJl����֎P*a��"�	�;�Ċ6���S|2�EP~�J�	K郮�\��P���`B��i�]�A�)	�.3�t�?3�Vq<Z�z<ՊK��K�2*�>"'\��tQ�)������y� �l�C�f���!۠�N�5+���lc�g%)Q"%�Y�	��\�!P��j��������&ib���y�)�pgL�ڹ��L�{ᯫiO�b�G'v*[�ȶ���:���	�OF��`2��Zl�j��<n+K����~��n�0X|�����;��y���Z%h+�X�w���n���H=�ޱk62H`���n缦���Yu��fJF�˿W��ȝ����=�eUj�Q׎g��@$�p�9�K�圠Jw�:۹W=MT����u��Z��o��	�*{�3��' �dl�c����J�+�X�>4�E�8v�.���D㹸��X`�X��,����yJp����he�#)�2�;���6�g	�n�>���4N��2X/~�s��d���_�k7��AP�rn�saQZc���j1��ծ�搏Y�YK7�7����KӾ��A�=�-��T����Z8I�?�W�K�_/��[6[�f[�]B4�cʏ����wa� y4�Mm{�x@t���B�4�v��۰��s;�4Y�ur_M��h����4�ݜ4��r eg���~v]�=���>�u��=&LC�f��W�<T5M��e�Y��P*���T�
�0�D���������8��]"�}F��7؟%\���Z��Tg��h��,D�N>��M�T�7J[c贘��% #� NA�ր��&P3s��2�6y���������/:3������޲8���j�����=�l��t
T�Yb���f�����=��>5:v�P�i�(Ȫ#p�;i���B�&���:v-��dN9�+BP�׊ep�ڈ�FR��T	��:21^kH�95Y�=s��v�h�bBe�K��Q�jl������8儓3��=W�*t	�M��|����6�y)ű�zrh$1��%G�k6��]X�u��
OXS�Qӳ��S�j�%I�+�/4��Z���^�_z
�����ʑ��B���R���k�;�Z9�U_r�Qe�$�N���*���Y��N�������xw�%V=-﫨�kW�뵠ܒ�$��4^�K�?�!�^�<74_��In;ġ�0�T$Y�9�Q�R#��D�,8�;<����P�\b9��E;����}�X�Q���G�D;���D�.׭�^�(#s�t�P��"�X�Ԫ����9���ֳ����)K�� ��ॡ��9�^� �#�R����F�|�S���sPx%_�w���mP�Z��8Vjg��J���Ϲ3x�h3�j��8e<NI��[��\���)nBx��F��NG���hH�c߃k^��ld�S�l�ńt��z:�J�"7Η���Ə�tiy�H�|єmf���6��I�C��>�`�|�4���36�/?����-���N,�\�~%�z��^J�e����P1����[HcU�W�N|LH������-���.[sk�����)|+w��p�B��{���b���!�`��ɔ�lRgI���{�ё2'C	��"��v`�f{x���yw���J�dw%"�_�G�x;��$���4uX�S�RT�S���B&���ś�����8	<p}���M�Np��e�B�M�&��B㶤�t�(�bг5온�[�s�d*�����t�4�ћ�V�7�Op:�C�J0>�2�J���{�V��o#���� g��5}�ala00>�[?\Vfab���\�G����& �-��k�Ry��x
! ͱ��٤�e�8��c�U?�p�u��	^����A��U!Փ(U�Oޤ�m1Z�o�e	�~�����1�o�^ ��s�'7�K�܈��j��)}�)r�{S#^6f�/a��Ʋ�����.k����)c;8F��"NԸ��_�$����1���8���cn.�*W�}�a8�wP����D�HJtK覍#��B+z��8a�;�[P��Jˉ�t1��ҧA�|9=D����7A�ǀ��+�]Ӻ���&bRB~�i����#��T��v�\��)�h�YD��
D�{�+������'(iI��!m�7t?ҽ�5���M�J�?%����p(���ӿT�c��%�l���w���O��K�tB)�ȇ`��C�_�A�n��MA�Kt<�C:n�n1�Ŏ��1�j�	]C '��4��C�Ơc�n��|i��EA�۶=f��e��#O��mE����0Nx�Ի��� c>��S|����S�$��_=x�Ni��ߜ��
֛�]�	 �l�'�E':;����ˤ��0��,�p��+^)���a?��==4�4�Hd�n`Da[�j�(��)�J��B�ld#��/���-��V�^{$�ݛ=�0/f����s>d���E�8�{�\�S>p�]�aX�=Z�'e��ܶ4;I�,��#�vP ��qM��;�x>I�ɺ`dK��v��م6�@�yjt /IH�i(��D�'sr�5G��c�&�vWQ�������� K��@@�B���+l�懺��S^���y�R������x��Rs"��FyHDZ�U�N�P&p�Ȫ��}O���"�m,��A=@���3j0~�t��s���C�?�*G&�Xh�׳~�p�_�Ŏ)7�R<��o��+��2J���Q��$[�@wq�uѡ�_28�|����\E-<@Vq���8�1��X�4e�D���km�̀.U&)��c�1"� ����a���+��L�J��Mi��ժ�^*�Z�:�� 5ڶ�jy3��J(<x�}��ĵx��v6\>�$�Y���Ƹ�F�~UH�Pj����}�GDϟ��d�6N�mB�ph)�m_r��P�N?����bg�'-\��p��,��zSP��VfDx��wpK,���I�ҭ�f`TA��)��8���� ?����Ąo����+�jm�[��H��Ms%���Yշ������
��ORЕMp�����Ex�u�ܗ�Is�bL����1��NG��;9���	{�(䐜"M��O�օ�M=�Y?�$���	���4�����,M��O�j����ʂ%r4~ ò6ړ�G��m"d&�c�7}����NO�<�@z����D(�~	.dK:���Qm�ѦF������=�]_ ��Wd�i7N Q��I�C�I$�����A�^��/l-8쮒�*��	�*�k�<AB�t��	prX�}{!��rwϫ���R��s�J/8m5v_�/���'���s�R�����1qZОt~.�V�m^�(y)���gF�ˊ������4=z��ھ{���;HV�Y�˙��\�-��(�'�p5y.�]��1 �R����ŪI�i�r@�af :��r�[�>��m�#h���Ł��]L�;�Fd){�V�<u��)��<��LO��sV>C�Y��h<12B\�?Ҹ@��;��Z���b����H��� ���0_HfJ��y}��K�"��^�1K`�z�_*��$∜Ƥ�Áf�mdYb�X��a�:D䥩e@�+����]A$8�� i�������6����������q-pp���|��J���H㼃�YV���~��`���E�im*z�z�߸J�0l��2@���5�P{a��Q&F�f>3cʄ�Ϩ�>7�9�<_�,�%2~�Hl�4���VyKiwF~�dݱV��ȴ+�y�yXh��� o�+�1w�2��T^��+������v@{u�xk֑ߜ!�B]�pm=q�50�i�['�ӄ{T�!��*��s\�֦>Y�Xb��}~&wX�-6'�;��f}?y��Fw"ѯdrˢ�[�BN�T��߂�?Ȃk��X��z�$�Al
@����q\'"�q��\t�ڼ�36�i��ZYl��
�ژ���qG���"#��z�-��i6�.��u%^2YU��3��_��2bܩ�k% {�mu�{aw;Щ�z���������փ8��ш|���6��q�̱��H�ꯋ�o�(�I��Tg�6uAuiʹ��[�����"C�h���I����(	��'K�������b�k�� r�>�)���[��Ff$[�mT���c����x�}�9�!+}�B��_�
\JY��������*�@�?Ga1�. t����1�)R�w
XF�+*5�sE�y����U��������c�r��s��P�:�.�AC��(����W�u����_��"Y��يA@MCB�E���/�zw���6Gm ��[�[�f*�鷋9�����E'8��ƭ	Y��͛w�}�}М�8L#?3س(�̅�F`S)���7�?�<�/�#����UP��d���q\Gۭ��Vn�z��D�;�w[����!� �C�	~o���X�����l��Ǌ�R��X�.��Û�I]�j�g1`�T�?؊�_%�+���F��!���6����#l�3Y��(n���r,�hM3�����5�V�s�)e�x�ax���ϴa>�Ƞ����-��Ԋ�-[<���2ǻ���]�L�$\��j<�~��Z�@�L��
����������Gɣ�A��Y�T�/�^�ס���G�i�A`dO��`��#��5J
�F4�oC��+z��H
r��!�d���dɞe0�������Tֱ��{��E��Ѓ�-��S�@�cU��#ٌ�63�t��°n
��5np𝢧��/|����.5��u���M8����0���N�a����E�[�@�[�+���p%�o?��-徎v&��13�`�2�v�r����'
��5m����綅@��0/��\�j;��a�ʷ7(���{�(�"��*�'������z��]$���#�Fh��_ ��aC+�>+R6��O��_��`�-de�P�H�B8�0����}F+9%�}.U����)���V�$w#H����)�h�P�95�!1L�?��?��vג�=�#�,֨�Z~���v(�:>7[��\�-�,�`5x�+,P�q��Gf�ܼ�,kZod�Ww�a��W�R�'��"sC�����cJOz�G��ɸadи�:�4��i��)�j{zS�n���8نR�q�^�p�!q��{��^h��II�Y�6���@ά�6tA�7q�L�(d�u�c25�m���aa����(�H�2�IҜ�5�g��Z:�>��9�ebL�A�����`!���p�_?�.A��uS�T�s�^"��ꕠ膷��[���	�w�yĆ� �Om�$f�잗�P���"�W���c�b�T����!�bO�V̫�NYKn�	����~Nd1z��h,� t�H�:�(=��������fhh?܇����I�a��(�Z��q����z�'(��OL���o#��IU��<La�
t������e�O�����]9��)�o#�#i�Ueg=ʨ�ʹ�.��N�V3cX�Zߝz"G�b+���Mk+�o[���8ؙ���sf���a��@eA"5̴����y' �ڰ_�y��G�NH��0I^)
��VK�L���O6���,Ǒ�y>=מ]�E���&{[�?�k&w�W�d��!JtD� ��e",i�����R*��^N�"Q�<�=��ծz��K��}�Y	��!�yc6� ��Fܫxj�����S��NM�4�l�{i�B�٩�E�����G�,���3�%�xe*����O���`��@�?l�i	��%^?����3��^U�[Ω��Xy	m�)���8�������J�*=7�b�{%''��V��(�����a�`�D��p��^�qC|��y8?`�dŷ4�DىrN�j���$��v�l��.w�N�.^0�l����{��N.F���+��7���+YS��</�p���)�"\�zM��#� ���ha@
D�����e��o�G��s	��V��@�!��t�=@	�IZ�A��<��XY��+��NE&|;��E�h�t/�����rL!���,�w�E�����f�UWT�9����C����I��#���L����p��zf�A~1��n���A������W�#�+�A@a���x�D"Ҝڀ+�� �����4����~h��|��wnhf&�tᵙ��k�]o�B����� ���K�C�`;Y�����%���r5ݪ%�Z{+�*^����3�}:�%���H��=m�(šL��W:S�d��sҶ�/�珲#_bN�ͼN/y5+b�Y��t;�����-��p1�a-8f���4��`����4^��_���ҪZ������7�4)l7v���`�s�Ɇq�C��lc�(���4�ݘ�u���ϡ��`�$�RY��0�����L-��O^��F~���#��b�L� ��%% m�O1���tu��O�0�(��)���]U��(��j繁T����E�ț��(��BѸ�2�U �����m�}]��{�"�y���L�LdRfg�f�o)-�!�d�i�$FZ�-؃l#� ��糁�!6����oE��5�kX���
���,�-��<� GqKA`���;S`K},���8z'f:�$Ys��gWէ��Y�Ut.��m�aM+=�}��`�S�ӟx[X��ܞ^Cf����/{�,��,h���$n/dt��^e2.�[������X"���ڶ,�ܩ�J'|�d�l")��[��4p��L�j��L]���e��ph𘙹1&:1�9��~�2<g,��j�����
����d\�AH�č�Pd�wPAs:�ȋo��Rj�P���g�tb�JT*�R_����X�g�@��A��ļ۾c'��x��<��X[����Ǒ=�Lu�$�ψ��s��
����Wx���eLk]^�#�ۡ�aC��Ҩ����X*%��ˤ���1�4����d'��v6m/q�~q�&B�8�<:���ϻP6i���ü[��Ώ����KdJj���շ�DYN�do��w�ￃ�~zZ'��������Z?O<F3�� Ff#���P����ʅ�gоW�e�o���a�ќ[����
~ҥ�)��k`g��$he�B*��o韷��a�l$R����9�g�mط��V���h�; ��snv�8�����cy�̊ �:dzW�=4;`����qcZ@�t��PÁ\��6
����&��)�;��N�+���4fI�eʳ�%���Z�����NՇ�o�+ⴑ)�����h��볳&�I��p�U���I_��1"PL���	�Ӡ9L
���1"�%T�d���G.���b�/W��uBۢ���k�F�� ���}�0ɇ����stt֑��:����VMK� ]Y֑��Iب��O�|߫ȋ{x�[5 �4��u/����89��;��mv�?��R.ȭ!:�/ ��F�"2G�@9I����z��L��0:*X��J{F�/K��)��M<�1�޶�CD��P^H�ܾ���7�9�0͉�6���W�D�o���|J�<�$ڲ�p��Aj|BF�d�g���@���#s>O9�q�}0����r�C��ew�dӋ�M�Dڑ9[y<�çs��cx� i j��wB���/^'�n����msiO!'��}w�'����Q"1Y�=p�́�w8���Ϫ8�f84r�ho�K8�y����e�ܦ/��_�Ɣ�o����sj�^���;%v%�����h^�\��b���%-ٺ,P��9W%�_
������Fj�~I�:ýc� ���J����27r�cU,kao��<F��Ɖ=���Ϯ:%�Di�*��f��H��B�5z�NF��������1���x�r�bV4x�@󭱿��I�rL�E�B|�� �I���>�ϕ��:4�!4m���Ig���(Րy.�L��
�cz�s� ��S�E��p�؅�4'�S��3	�;ϰ���jͼ���˷
�#<�'yv�q;���s]�U����]��$:��4i����i�������K/Q�"_�aXI��RT@OHc:��F����wa� �q�Q��C�1W�d%��6��;�gEPm��Cn�Q返��"���"̷;�[O��C|�`��5ˠ��Z��yD:�M��eſĺw��6��[Y
��}7����o�W``U��.��Y	�:%� j�3�������O㧶�.4�0?�����>�{�n�R��ʲ�9�~?��"��ցʯ	�l��{
����_�u��23?;1hC�&\�� GX�)�: C�錻������!�wpg�Y������<vq�i�"�`��j�}wf�,�Jum^�&�H�^��.�lDK�Ԁ݉$w�t�����K�pb��gn%-�٫�q)�;^�\l bƍ'�s��� ��<Ål%��
��L�#N-����0���!�# ,���Ԍ�C���^���n+����m�N��HH���xC�Z�2��2��h�k�>O\_#���5���͘�)�D���q�\Z�e����q�2k���o�O:��.qc1�2LoOčk�(Y����w��\�T�[����:aK��ޏ�ɼ]��4�6�(��_��Z�*g�0@�2y�7���u�t�7����.�����D���=޳}�K�% k�z���]�uX���ǟZR<R��u!�c��ok�OT4�#X4*��ˤm����ܽ����(7H�����G$����u+�W����z�gU�����]��G��蟀ܳp��P\G�=J�N����&n?3�o�3缇��i����Q���͞5i�b���(�x��(��	��B|U���T�4`�X��1q3lKq�u4\Ӏ�f�\8�XmMM��`�f���D�8s����3�p��6t���SU	��Cl��ty͊(�q2GB8�K �YH�OMlw�e�2�guf4i��h=\�S�J�/E��L���J�RG0�URK(���O�P��Xi.1`�`J��}}�����+kJ�bI�~��t|`E�'Ϧ���l���e��bJGd�䡃���=OD�!U��w�v% e�+t.���<��{��pvL��x��x��Pw
�BH����=u�p� �<�m�sُw��f`�.�����x[= k�a�Uj�x�O��r*ċ6YL��15y�U�\5�������9���A�� B�,��hH����0e�(XA�N�1O�>�B15��n4{��K�F�Uv�@Hf��'3��P���<��Jz@���e�x��Q?Wٮ�Q[:M��0�<OwL��6ҁ����+C缦[�r�gC;�4�u;�ÿ���F����mc���<�R8r�ALGn��F��ud>ɣЂdY�l��!�'��G�ڐۼ1�U���K,�Ptl�M�^��[�w�~pCL������UV�MQ'(q���o�H�����Ni�4_|�F��z_��:�q~�[��R-*I�x��R�Zd����?����>��,e�,9Ѡ�J��7�!��=���h* q�4χ�K� gT%����K
��C������Ѵ/����N�S��Vziv�Å��^!�_�{�eP�k���(�;���;�7��ħ��џ�R��9D�
�6�&j��BXvUD�Mh��9�/��a��X��Y�t���� �����m�' ���oL�@����>��YE�lɢ7K�ZAt�葒�?2��{w�R< ��Xi��wG�c��������J �`~��z�U�"��c[�� ����Y$9~q�NY�Zӌ��,��œ:�Ý�*�	�е����zv��:��A����di��t�?�Lb�N(�0�ITC:�ޣe����EX��W�u�ciX�%��wL#%�*&*6�wD�N�+�t��*\��l�Ǿ��5��)AZD�@���J�v`�0��0Xk~�����_ߌ�����躞�ϐ��w� �<���bʒ<�ɴ
��1���{���8�6օEt���?c�����\���y��*�|KrA{>H5}��+E�)S><�gy-�GA�3�$M��#��ۦ�I�YTg)xGj����<�F@x2p痵y6�xcUˀŖJ��h���@�1�:�@�y�o㥭��k����^��|7��L{�H3��|F�|�����Iv�7û�M���s��>窥V��,*���ָ}SR(�? 	��#.���uc;T�p��z�f��F�J��&4 \�<lӊ��]'J#�.Y�~@n�%�w���F�L�'Fy{Ш�u��m}1�j����kA�1,B�ː������X_�p�q����mOv<|;3����@�8����w�fUY�����Ow�c�"Y�9�}S^l_�/�5���SS��K����Ҥ��GLؘj�|i�A���ݎ�����|w2��3o<u�>���P�������vqd*{"�3��^��٠T��t�d�|��[@��9��e�ޤ��/h�;F?@����Mb�|2lu{�
{:��>2�1�7�N�������R �g�^<�y�ڪl�n!�f&o��to^�� Gѽ\5��/��*����s�fh�5i�Ѿh������yȧ@y�������#߳^!�L�k�sEA�~(|��E��Kp�O;٠i��bd��X�N����68����~�|xA��5তmJ�XT��wd��n��� ��#���!F��W��)�?�����Z�W�i��{�P�
 ��R؀8_K���7�Lyf\M���)+��`p���v�Ы�O )/����QW��4	�\�=�
�`�E������P�����"K��e8%]�*%՝M��.Lv��|��8�W�� ��kѰw��ȦE)�;�>1��p+���<�(y�dL^W[33��B	���Z��t����4�Ե�6륲tc�駨*̡D��gW���F��E߶��B{��l��#��[���@���'LŹٔP�o(5���:��g�%YV�L }�� ��m������YZl�4d�p+z���|�:�4[/J�81LG�_\B��z�{����}B�� �1'o��d_��1��֗[��R���mΑ�U��L��BO�G?�-�����s�W��Q}�V�R��˄�:v=��	d�5 8	�LSa ,���o� ��������aw��f� Z#��q����0�j�߱weVdl�975S���e?z���.�`Y�3��:~��Vr�e;l(7�m����O��W ���.EP��U?���:��� ��}j����#�F��!�~�3æ.�&>u�k�B�p�*Ɖ�?@�,��]Z�Э�9�!ʂv�z	���W�pb���E���my6�\ij(/^�;��{k�1�=�ϴ�Vb�<�ҷ7e�,��^)�-�W�ޓ]��Y,[_Ju�n���OX�>��ޣK����Nd��"��A�l�_��gV��P��¢n�"�L`\��i��������6��s;�I�1����Y���l�P�co
4�}��p��9=�)K ��T]X~�e\@��;w; R�1���i's�ri��	ɖޯ�ͿJNI���Tv~svV���Ce쀷�9�;��j�3����S43�����]��J�w$.�[[j�-��'6=��U,k��|3�^ӖYw)^zd<W;���pJq�n����'r���]���A(cf7�4�#u?e����:l���[�����T*]��weY -^�rF�/�w$)g��+{� �/Ē/����y�x
�Z:C�}��X�z�&˙��)]�q:5{�Ȉ,z[�&姹I����^���M��U/�'	��S�+v��-H�V5��^|#���L�mz�{ �Ŋi��:�жg�Z�-Ë N6�m�/*�d&�W�WKP�N�?��漢�ӝ�&v������Si ������q�m��d�x��D ���Th'��(��Z(���ǎ��Emm�j�����n;m���ÔY�{�NY�Ӌ�>��-���wH���o��c� ��K�۴I�t���w\.���%��R6%�>T��~I&�Ϻ��3%I����i�ܰ6������G�k�� |?$�E���\%!�>��+�7x���"0�Q{ z�C�޼�O@:&�-(���]9�lq�_:��K�]o�X(r�OBj-u5�u�"�������I)MJ@�=�;e�e� ����U��6�M
�������ٹ�0fHVm(������cj����f!���E�2r<< Ih������W�Gr>���r}ݔ�>�2����ü`��-$n�å?�t���}~��ٳv����xB5��8��Y�g��@��*h�[�9���1���Bt�e@_�6��ɴ1�U����/{� �^�g���j�*'�X����_�XJ�]�r$ۂr��p<x��3�����D㰧;K��gر�`���<�_E�R�Z6=`b�r��� ;��CQ6��,,!�hP�TX˸0�ͭ�V!�����L���<�R� ��J3�yw ­c����uZ2����j��-f��A��� %ѱDTȪ��Zy�B���0����g���T�Z׍�ۑH��Vd�1�܈bc���$޵��+a���"���K����j�y��r`������K Z�RQ w`�A��e�Nk�w}�����*C�LJ��(ȎKH/I��Z[��ׂ����޴D	�� ����K&f{H�I����8&G �cN�r�8c̾��%�<���90/:��s���2���w��Nl������	�8 {�z<U7%����B��W�A��hGWR'���y>�����d͎
a�ha�L����T�S������j�H`*�K�Ӏs�<Skp�a~��q�ۜ�0���3��ټd���m*��m	��7��Q�P���]��E�Zzxj��<v[���G��e&��Wׁ�=��i,W��e+��|���O
�$}1[�PEtR#O-��:,S����=>g�Dd�xk�2���.ݲ�ҽI\�$�su�]�0��0U�����4���hS��nK~�YB&��U�PeA���q~���ݟ��xsSE�dm$ٴ�����vT�=�!%c�`3�3䭕�g���Z��IU�=CNbvE�S���nT ������Z}�$]ʥ�,�L�xļ�¾�0vݫ���62���8MפZ������]Fa�D����Gg�������8��TK� x*^���KD���w6�P��!=8f�~9ΜE�m��5瓝�:N.g���ɆIF����J�X,j���^G��;7��* |8�?PQ�VO���'�H��A|��p*N��IQ�tAp�3��x��b;�叿=x
 �Eڡ�rY�)Y�k踻�L`����5������9�:�=���-ֺ=s�>�d���&�D<���1?����^����dh[dN1�Ɂ�n�n�:ZހT�����R��ϗh%E۽���ʍr�*���� 3V��.�J,�_�5���OI\�)�U�+@0K9���rѿ-Y��ƻ+�`��x����
R��+&�zX�v����Jk������/��{�l2��zg�K.���t���7�!���K�Ȥ6�7�7R�������<#[��f�\�ʎ	r~�35Z]�&#��2U�����&�7=��ʧ��mo�ǚ����j�� �?s[l,�c��lw��`e���a�e��P��;�� )��鄅���P�Q@�gL���4��=J��� |����󂒔 �;�w�Y~v4�5G�mX ։��	�m������J��5�;��0i��_d��o��X�a����S�3���/>e�l�T#
�������V�Tf%kc���0N���v���)ɓ�a��S�����|I��5��+��+��+s����/��16���fd|����S>]��s���"�J����C���GmS�;��hϡ6C�B>�D䧋�@�	m��̀�@�#F�9������L.�c���4�{0˔��s?�f�h��ݷ�=��/�B[�[2B�Y��̠�{ ��L�[�鄕؆��[5z.N��%�>\G����g=д^;$�-�y�VLL�|AgC)pUƸ�� �2��Q߹�?�V����ATLp��U�4xyyd=�#����J~Pj�ŗ�:��
�kl(�Wm���kg..J�U$ύ"�Z��%6Ny� '�����i6��w���
�+�1��.����Ƽ�6�oS
�_�ɕ����̭XM�g*��v61��S<���J�a����Jy�v�Q�#�I�V�wc=B@Z��:���Fߢ���ϑ�I�ʪ��H�p�{Sg�K]���	��*CxLaM�=,�D��2Q}��4=\������!Ϝ;v)M2���e:��{��_������N9+�"�4u$�f�N͢:UZ�7p��F�z
ɠ��t$L^[���5�������I�%O7T_�����Q���1J�-�\�g�jM@)�������Fl���J����ٗq�Ƨ���+ӄ���!ӗz|�1��q�/ٱ��9 W�+��:(�y<v�����O9����u!o�x=�;iksyr������dMӺ������B��I�E��z>�+	Ux���g�����@��\y����ά�sM��mB0�P'�f�j���h���0���6�R!�����>l�y��Jg+�[~���<6Ik�c�m� =��(���:+�8����y&٩��Л���� zc��nVX�
1�E�20.�p; P�R�a;��s��E�TB޷����y������;��alG�mnN}4�7&���®���?<�	�Lv�d3Z}o@�t�e�����`%�R,��)��+�c26͘n졜�?�̏��d�����)�}���ҫ���*��0WZ �0o7���*^F�5������!d/N��:>\���O��^��I!G�[뵃����-?����F��rp�����^ok�.8��*D�h�z��{�=��=%wF}���ZR�m�пV&�nc�Cl�v��S�Zx�x�{�h��
n5��4˼��Jk\D� �ė�t{���?�cbh���:�d�
Q]P��\ګ0�j���~�T_v��8�e`�fF�����w�p���ʉ����D�w~��0O(�l������p��[ީE�d���_w�W?��;�O��<�Bi���W2k	�)a1~ڭ2q��qg*�|h*
)�-4W`��	󒎓F-�@�$+���A�ӽ�.?����2��9<��V��u��7���16���iLÃ@�ֺ͏y�s.͇D�ͥ������_�$�b���k�ڗ�Rn��A�x��	sq/.?^k�`5iu=;+frF���W�-��ఊ�V/�]�G������s %t)G)��H(���:�d��y>�i��=û?��[��m?�E�w���zݙ|���E�Cs)4)`�pI�=	eBo�+򥩆Μ��m���d�t<�/ǂ�>���kϜ����;��T�+yN��_v��e�-�
�Q}6r��%����`��YX���ƿO��J�N�o��[zP��?��Qs�6M�Q��eJ[mF8�t�h�(��� ?��J�&6p��@X��|�����(�vt�̃B
�ɢwW�&/����!Ԡ�=��U���C����4��+�I��Y��f�5}�<�'���edT�L9f��ޝ�}�E��+2���Ry艘+O���|(�a�T6A:/�%g����U`�|Ń��l���j��֮E��SӵUX0y��A�ݒ��E����V`�
ó�N���|Hy(���4��҂���9	��@r������ ;��U�LR:	��T���sM� �-5�/Ӯ����\��Y	���h�P����{i<���vZ
�t��"2�hQ�]��_W��I%/���a� .�&�2�܏j��yd�Ի��/V{�e2���6����o��nO���К�n|]���~Φ0V�&NQ���Om�J0�a
��";w�B��ޚZ����z�$�u��,�� |����rA�,�HO}jK�~P���L8��s�<5%�@������`<�nG��X ��2^6�j���]L�|l�&o����� �	��)�Nf�vMa��ݰ�W�Iց��]϶����oV�I8��t���������:>r��y��9+��
N\�۟D/7��
�v����s8����{a�x�@�:�H �uD+�i$2�ɺ�{�*�?��}��u���͟�Ȑ������
��z�Գx�h�r��~9u�&2�:�p<?�X�£�v����[lJ��{N�z�v)��,���?(�e�+'�(�e�跮FЈ"G6@K/����_J1����;��M�'^n�֡6���>t�9�8n &�`��ӳL-��}*6�.�.�"-�٤��/M��<�\���M
�,���=2+���W�}tM<~:�KO[.s�ۯ�J? �y,^�A��;=��	m��N�в6�=��Z�r����U����b)�E��t��rg3����w���4�H�l8�ؗo .D�bk೴]%�0m��~{\W��W���,n5��@,�g�\xuI�<���ϯ��W[�������r�/�$}�=QF2P���s8���=i�E;��_hµ���<:�>f���8��\ޱ�GƮ��9���)RA��^UON�$�R�R���/���g���5aB��bz&)���ٺP	Fb��
ݠBx��=���m�V^�n'�����އ�-���G���u2�k7�����6d��+�vg����QDY�[P��|m�0�2�7���/H�C�[�9�I�%8�m2�����:�:)ǡު�W�
�q��
�^� � ���!v���r�Ԭ�)�4�1����IG���\�~� oq�{�ԐD��/��z��*y�g5���s�M��[,B�)�_�Uq�J���:[YS��Yn���(�`N͖���h/kq�"�Q���ly���nە8�AGu���e(%GYv����$����?'A���ح�ݱ�C��5N%'P�]�&� �W9W{k�`�ܯ�w�se�@��a�fz�M�ʶg�U��/�%Gۘ�^N����j��4�|�o�ׁ��y�
�b�)�q7w%�H�XI&]��m��1
m�ԾR���F�p2��V��mU�{�:'w�m�9s�mOs9�q��E,�d���m!)l#������Z���,���y�.�_y#�7F��ix�J5��
�<M��x�������y��AW{M��(E	8ֻWF9c�m�;[e��g}�ɵo�Tp�rGl��a�#:�f�[��g��v��z����}���l��1�Sw��0Ɠ�v/Ԭr��#u�:�?��r]��3u��'�7~��G`��3�U8ɢ +7�'!�w�E�S��%]�XӉ����v�.�w���i���1�=�p��w!�5� e�l��ޥ�-`�s���"���Oa��#�� N�
�9�Y!C�d��@�P�Bל�"o��>�q?��a�i�}C�F�+nt�j���y���Èj&�f�!�|�K���c��Q}���'j��{JZ�5�gc�8-V/�s*�Ce�x�+|/�z�|�׍�1\�'�_�}���-��>�3?<�Ѯ���\��5O]B��=f��K)5��+��B��r'�:ңz������U)l짰_K{1�T~lgw�v����~�8S3+��ҥ�1����%�k#I�#0��,�9S�)���mS&�S5f�'�@GmJ����sm�D��Ø�k�f�
�N-��	خ������+c�tN�PR� J�0��UrR����oR�I��e�m<����y�)� ���Z!I��?�3	A���C���������y��j5kw��)�7]���BgS����01Z��:^V	�Q:k9$w6B$�{��֊U?רr`[2D��sͽW��j�do��%��_���C�||�MFl�EB���n�\	���Z8BM'�?�9~RI9qSLˎ�:Y���U�a��R%��ޚ�=������&��,�^�]3&�jwG��#F���DFނ�÷4;׍;s�TZ^�[�����ûȯ����Y�&������E��,��ڎ�#��%@VoY���V?�f����0�8���?�����~os�v6>}z�(�N�'�KT�Zn9��	�7���}��,��q.��16ǢQ�_>o�9`�$MK+��̷L��V�wX�V@�,oAY(ؗ�2c��o���	I*)j
E�	<�Ә�Z9{�k�RF'� mU >lta���u!-��{ۨ���Л��RAGyD����	N��@�X�߮M�����Bx�Y�d��넂5{��#�7㺒m�<1�#9�\�$e�H�T#���[#��ȱjA��{9Y������ߒI�P[AY����BD�!~xx�m/��7��ᅎ]�*�l/����t�Gief�3G9tP�����Q�S��`Lq��2����`&���asꁔp�0:֏;�{
X�i�7{ ���Є<�
Xj� 		�&�|>)�H�r�d=6yN�b!j^��Q�|�N%zO]9��%Ŭ�d\$e��6�1��Guj�M
�Z:`���p,����:�Z��2⧪��N֨��aD�ҹ��,�f�m��E�ڐ���D�*�5����jT�����yTh����I>�mW�$����x<��g�?%����%�f��n<��Az�y1?GVq�ɝV�罶;�f$V��n�(~tF�B�������M8�9:\(�ª�L(���|/���	u�s-_,��8j�q�)��Xq�%�z\�1��ZA$��{�`ý�*_�̾�Dk���I�\>�5E��נ�	�8v[��'���5@QpE؆wZz��QO������9hv�{�1r�Ik[��A�i�\��E�������E^��\�-pZk�Y�a�;}=(��*Y�OY^�Z�~*3����/��|i�"$F`ULhb�]�ո2�d�-�Gx���j1�]�ګ�Ʉfz	�'
L�E,�"i�����G
�2q�+EŐ�i��\Q��@�h�E�������f0��j��ŕ���\�Eu���y�A���r�V��ت�`���J�̂"'�<1.���{L\���4!gH0E���u��Aq:��Z�_���Y��2��Nu����:O���p��f���z�p��hW�)���kR+�����ػMS0Ϻ�<��L��>�$-�%fz�Q�#�ΐ<�/(yNy�)���gF��^��-�$x����vp;&��j檬�3"g"�Ɠ��t6�Ɗ&YJ�2H��Jw�L�,9���'W��+ὩJ�oC��ܱ5+{P
��ǐ���d4f���(V}�q�eN���	;��?��T�d��T��H2'o�2�j���E��L���g��s�0K�+���D��\�.]��ħOp��zr�X��yj�A��!VN'W�� �Σ�������AK�}/�bZG�P�4�mH�q�`�<���"Gأ�g��X�@no��W��6�2	�*���֗�v'�� ��,4ԪK��� 2Vߔ�TI�Bߌ�--M� ���>q�v�zC=<sm���?1U�����<�?����c����J�lǝ�|i耇ӻ½l�&-(!�Y3�ni�~?�0h��}ؙ�}����Sܧ�L�Ft��k5����9Q���E���.pXZ�Ȁ;��6�Lأ�*���������G������@!��?o��F�t71�)/pȞ�q�|M`<ҟ}O�"�E{�%e}R�s�^�]Ujٝ8��7#m���;���s	��@�����?�5�!��}<�e�Ǫ��/{ug)5/3��ub_E����r��l嫬�Њ���)���/��v|�1IcoX������hS�3,&H���)���e��6���-#�M�y'ώ�`0�<�?���"�U/Ҩǳ���/��mo�A��8�<���ýBM��a��%z�U|ڀ��	`�ڙ��\���nD��Z�'� ���=_K��t�"��A��lYc}���@�Ht���Q�!�����͝ceM��<}��S�+Nq*�t���U�K��D �ܘ-�؟Y���/�%���.hDg�\�� ���W;o�x׹Ⱥ��16%<0�w���ɝ�xlmS���JM8�C��(�����ؐ�Ƿ/X�|��$}�l�TՆ*�$���x;Q��8��P��w|5#��tE�t@>!���C����"�_�ӏ�5���P�v�{��PYkA�CQ��k��`�рRu�Y-8p&ՠ-�v7+��hb���~ ZBÚv�gJ:�����,�x�>m���� ����"��P1�p��j����������f�~	�,RVO��e��t^b5��:MlAV���񬮶x$����Ѯؚ��i[m�3��O��`A}��5���8��)��~��(�+C���V_{>2Lߺݧ�2'�;_�$Z�r6���π�ȀQ*5���F>T�C额����Ҽ�j�W�)��|�[����=�vJ�L��pCwRS�)>� o�o���i�	А#��B|�����돬�;�)N��O���(�}"��w&��IE�R1������;�`�g������%��,���D�x�A��Gn��z�@q�'<-�J����z��
S{�RF�]~磈E���kʚUbx��x�9R����|��;̷/��BbF~s������o��C-�����8-3�O��(�$Ce�T���!2e"�@i�Z�$Ӝ"l)���������EK��=K��(r:���s�~��漫��#q!F��([�D&��/l�\W�����Et�m�S��He�b�x?\W_P��3���t2p#�U����	��D/��<2|Y�?���<n��D\��BJ��R��ַ�����Y:m2�@��{z{�W����y��$�T�Y���`\��m��"�Y���XF;$֩���:�˺��9��C�~����X吐[[���ѓ0����z7��)�~z)�UQ��>����}����/d���"���Վ%s8O�)[Ab_�pW�G������G1g(�vz�KjOT��1�g�����<*�Fщ�^��Q�-��Ԁa��n���f;4���,�xy���+𯛃Y�Qg깥-�L#!�+h�4' ��5w�X� ��dし�<3:�F�z3��b�l�?�BQ�jG�B͔��s���͘�^�"��
�~%A���%U@�ۓ˞�ӕ��B�
�A
����:�:ʴ��ܬ$�8���|mTD��n��𗞕�ͪr�dם g�ORy����?h���S�@�p�pp��c�zh0j=1�]���\�<%�Y�o5�r�F�	��ϱz�S��8)�ũ�T%:ؘ�䖦��όRދ�`��� ��0��Z���so��4�ײY�29�s_����U��@~�X}t)�v�~���^1��/V�3}j@�F��B�W�\L���ڼ8<^Y`�p%%d8�q��C� Z��������0{�/0y$��aj?�_Rj&�x']�B`2��cm �vR:	�$�qN�~85�*�-����B���C�Yf�M��1�[����q#���H�Kֱ-���l���M`$E�6HOk�������/��O���8�=�1�[$�Y�,p�3�����]|��?�pA*]��9p^�ď�1ڎ�td��0�J�k<͒�Xc/�h"�k6�s��p�~�8�yW7��В-	�,"+;/���*GIo��aOIꟺxm��*����j�Y��� �<�H7$	�o&�kQS�m�-��_��4@�M礑/PnDq��a��ňՎ�Ϛ�M�"��H���[I�I������>�Ԅu�^�wK1I��=��_	�9F��J�(���HO�+W�D����o�U�l�k�nn�Α$�␫G�](P�Y���\r�ͿH�f�a�!����8���!;zɁ���6�-o�n('�k�sd�Ų�J�|c*��钉 ������R�򘝘C��6U�U�U�m��8<�{��w~�j�z#�i�9�ҲX�d"!n��qVw���q{�����*l6N����AR;���b��\�f���!�XUE�痘�ַn�J���&�S?'�=�O'FhBa�!�X��k�IgwC84��8���x��v=ˆ�VX4d�b�|s겇��M�^q$OF�W��Î-Ҵ�h�Os�2:ɈZ{5+��eNf��N���
�I�B�:��}Q-4h���`�S��)nz�:3�%Hd3�����<�B�0��2�Aɉ���w&R�K|k�'J�_��bw=@L��)��o������ߠ_2�YԱ�Y�Z�����Ȭt�卌�Tޱ��.UeYE�LК�	���s�k�H'@�a��-�9�k�(x*�b�H뾇�vAީ(�Q�9�+��r�8��`�}��_�$Š$��1���37�L�����9ML�+�%^O�Ofށgzo��e��q��p6�ݔˏ>��d�.]�[�5���l����ρq�f��N�����N,�wA�(sXʳpa�>��Xk������g0D�M�.V���x�չy����{�(v�S�8��0�&8�cdթ�+]�L9�<N8��ޝ�����$ŷG���@�ܢ��_��s������v!U��
�Rl�'�'�!-�G2�9�L���;
0�t�ebS�歏��{�5HS���n�6du<1�����{�Sb{�|}e��~��W+�6�^��M���.�>!�9�P�K�c��\��Ҷ�QAs������@��Ԃ��}�b)4�^X~�Ǯ��c��X���4�
g?n�E�����]n�^n���X�8l��L�*&�S�֐ @n0�]��%��������M�T*��o�#�F�|J��CWraX�â����-�3RmD"��-r
�����ui��eg�[x���T*cIc����\ڏzi�	�,�I�tf�yh ���ڽ].�/�zP�ނ��Xu�O'��9@�H,u=g�����;I�_9�-H�N����P2_E�XK�O!�����(j����݂A���?�˛F�	ޛ=�8�&�ir�+@l�_��vʐ�p���Na��n�͏�(��X'sM�����atޥ�qA���H���-}]�)�ɏfDاY�����[��jI����_�:y`��/�h#���g4+�W3����dk�9x�"�����d���r��ZG1!� �`�WBCX�ٸD�L����Ӛ��C������ד��o�lULӼ�~���$ЖՔ��r� �g8�I�rn���H>��Pv>R��Ჟ�����`ɻ��� �:�!j�z5�� �?"ΐF�DL3�>�Jhg���3�� ��}��ئ�5�s���=R���#�o	[����+� |�S�,[)7g������4�>�I���yn
ee�e���7MMu�*ƫE���4Sc�rPA�Pm���29�|��!u��:��}bޮ�f<�^��W	SŅ㑘�1�6/z��E�_�Ȋܠ(E��s�e�ܱc,,������>H���k�\��C�>��%��U:�zj�q=��&rRH�j��z�!*iQ������5��Y�F0� ����ԟը���#\��B�p�1��u��nv<�H<Bct'rC�a�����~��d_�4K��}�¾�F?{��-���W��l�ҵ�snB���`[K�!�!V9��������[�'��3dmȧ��_�9zXv"0��������W#o*AዑC����k�Z��X"�m�<����A.���R*��HW�>f�
C�k�O�3r�	��+���j�	�A^J檱�_���/LFz8���&iyWg�>>aSY��#�	Jέ{Qc�,����	U#ť'e��OgE=��:2��h�:�_�NqB"U�1+�0#�����O���%.q1��o�QrDM)4�e�H�0#�a]k������GO��-�/��j����Յ�22�RC��%�d��c2=�T>�"_��ID�����4$�p ��:�Ae��Q�00$�s�,�9@�mf%^aK�tLbnEhl��٧�! ��C��>�U���z�4������l�7c�G��ri�{h�8�'ON�+k��m0�����ό�=8,4ug	�������Cw��Vs���O�ID6�*F���$���Y�����x�ok����/Q�Q��d$���v�|`��g�p��#A'm��b�g鍦��G=Jo��ɍ|�؁��z������ّV �; �V7-�B�%�԰��[@G��Of���wp��ݹ��? ���)��@��h�ƒ��ܦ#��c_��U���óE������s������K��G,*�q�K_"��	�GK�8�i 9��wa���w!�}XPr�3�B<++��Z��
g�p{ؿ�P�j���+�~3���7O�M.P��6����3R����B׀�EE�v�6֮28P�Δ3�k���W�#�DB�b�~f/У`%��8(_��#��U�H��6���o��[X��Q"�K���h���DG�"=%n��UO���M��gX�LTl5`����qrŕ��,��������>�e��Y�ώ����V��*5�����?����&����pL4�*^~�x�O�J�U�n�4Ȗ���A(^S���� >(�p�j%�.���֭Ξ��uĔWr�����r5�VT�s3��1�"��S:�'���"�?��K��9և�`&�0pa�u��ۻS:����<�=h��!*��zݏ@�m�H*�(y�x+k��}a�Z;��X1�8�^2��>�������Hw@�i��?�ЙD�g��oZk'��e탂���m�O ��<�Sj�	�R\�`�D�	ԷV'�Dt��9m�W�a�i2����薖gӟ��EDͳY
�1U����s��U�bg�UW�=#��:��U���mI��$ڕ5�i�P�)C����Q�V�^,5o�p��ʕa٥���y:�\��X��	g5�@E����dD�rWa2G�q2�&*X#13��OV����r%Y���!�`���4�iu�c���!�	�L��Y��-��$A�,�r��ѱ=Bv1���u ���p5V��6���]��`q4���/T�+>��o�emzrq�̓Z�<��R��^�J��36��L���f[��[�.v��ݳ�=�b��p���������P����:�@����o��B�,�h���9�OP�΅'��ܷf��~WLHof:ey0��@�CI���������Ϩ�	�a^���7��ȳr�y)]��yd��-o�8�1�rΈ��F6�;�߃�H	���~6������m���e�)@�8��L��&ˬN���[a�w�!L�x�`:F�̨E�����~/��j�g��d���?a3mh�S��`o���s|]V+�;D��:,\H��UA��Ae�c����L�4��_�v�\Jkڮ�V��+�厤������Ω���@�K���R!��������~� ~���;���b4i��r���'�/�����vSUD0�m�[δ,���~A�Ԛ��Gy+�J��ڸ���!f����2���/���r��r�J	�.tej��LB	x�baCV	N8�0 d�mf��(�x�w_%�Nb�_��.懎�$9o�1!؜����X�J[�zD���e>�~x��&�7	N���Rn���c��C���Vɒ�p���o����IUUߢ�� $O�"9���fA��!�\�PT��#��z9u�B��.*VL��ʟ�.��������vl�˒��?˲�m�W����W�ӻ�^ʙ��f>(;ֿ���*��߾�R�6C�������^q���s��)޽�+��Ƿ=%��<&Asp3EU}@S�DFp� ���*ME*�઩���@1�O~pǾ�LUݷ����w�?�]�v�R��A�2�>{W�Js�T��X�'>��TI��m*����j6�dO����T-]ɧT&9���(咐~��^;6� �c�J�H�q��Ԟ�̫��hg��k�z�88? �pk��f _����Բ �7�6���)�#V�;���e�m�Yx��������,����;{1՟��Y���j�����ѿ��5I��ң
7�,Վj� *�#�f��?������3����s����Lޟ��dfx���K��(�X�v�R��kʻ���7�D�WU�_�P$��:6����%b| 4�m¨���l��5|`��bò���g�Ԯ��&]�_�#������t�*�H���KHMO⚜-+_)�B��k�3�R�M����OUֹ	����_�"�����5�j��_����4���)�e�>G�P��qP�ߣͩ��tS7���\c`�q2���Z����j��[��N��K�}��пW�nkK�p�^�� ���M(��wA>���U�t2��&��#�u��@ẵ�B |�f�}�P���x����+��,��c��Wx^s�<��hzO�䯨i��9f�o:�rag�Ҕ������?y�H�xݞ�&���w�Lqqĸd�I����R��<�&R՟v��BjL��mp��~ߟ�7瀲������s<������[��0L,�3�CmM-BZ�{�g#���CW�9�Av�c��^^ �����{1���2|�?���b�3���u@���7N,"�B��O!����J^�r�Y3�xi �ӱ=�k��S��BR�/f`��w���I���}���U�l������V�{��d�>�J���٪�I"Kf�7id������6νmԮ����KQ�x�iCTVA�pXE=��H��I�����"�"W=dxʹ��"��p�cޣQ�?��״!�.x0VG�+�B��n�'��Q21���y+Sa�WJ����[zc)eMd�k�p`��A�`�|��"[���3] "n��Qz����#2^�<u�%s�{D��Ԓ��n:dd�
�i>�<� o�B��@B�M�-dIP}�gb�qA']̌���z����'JP�<[!��Jl9� 9�4(��z]4��p܉�GS���al����x�N������F\���QY��ڃ��Yj�����	��??�ʺQ0��ӎcJ��S�m�dxG�������3S]��u+��X���\�6 \kr��~�_��~暏�-@Rݏî�0s*�~��pz�^DE�3l��9��5�B,�'eq)�T�Y���Z%�I�@�r��=����L���0�Q���
����pq���\��*m<yZ�F���n���6����i�zj�'�[@��"j���=�1�Nw��8�\�q-�,Q5�Hh93��5n�J�����4���F�X�h�MB����XT���֦f%��M&N`� �,�b�g��@�sr��"D��|DÛOc�˗�M���М֫�\|*�3!7��m���0=���p4��8-�� m]�#�%�t�O��2$��N�:���~�R��B�S%��S�%v�Ǥ4\2��_�������u���FR"��+,f�7��`�A��u��cj��Vk���	�-)P	����Q�dê��Hϐ����'&%�^a�'>ِI��w��1	� ���ْ�xE�:��J�R�R�\3���?��	�	���W���B��p^1>g9������s�^��7d�e�Nv̴5�DK�M����u�/�4�����~����,��Y��i}�<��ⶎ�粍����d�)͘Pe{���A���=Ҹ�57uM�s�«���a#�P�h�A'�I��$��UX���4���?��Mk�ځ���a6�8���͒l�\)�&��������{樂�c���su �*\�9�u�O"�v�U��DP�r�=q�ү���x��$ܒG�/܃��
u=�����S����0��H�Z(�}Kl�M}�I�O�y裑�ݐ�y���9.�`٤�p���j�8�b]��r�[=1c���������Ȗ\�[��q�lGʵG�1�b�X�}��+��W���V
iFN�Bp��}��J�K�[0^79vA�1ym�M[L�G�l�`�៖�'rtS��|N?�W�~rQ�8�P�ڧ/[��/��=�<t���⽑��֘?�zD�~3�ă^.��r�V��@�z���7dWr�w�i���Ϛ��C��2�t~�J���&���ZͿB� 3����X�=���}�����vV[h��ߒ�-"���*��(�N�"��2��rA��HH�z
rn��q_��2|�t�����I�_f�5��,I���5Ձ���_ɧ��x���#WY��C\����5	�,?��GE
�LA��a��@m<�4�`$� I�Dej=>���B���$����H?Q,��p-X����U0M`i�
�]����K�D��N�����3�:t�Tm(r2�'?$',>�&�Ź�P�����qE�K`({�S9	eEPo�w�� 3�������`M=�]�Vv�5�U>E���!�/���v]f����ƍw6�"վ�KNO���4eK_�Bڤ[�����F�3@7Q:��y�!�W�`��4}q�b�5�"bGO��u��2(�>:����'���J��~&F�Ͳ�2+S�uD�߁��ۆ	G���h����e�\�A������a5hc�8����hZaq��[tv;��$>\QuW��m��QH򢰭�,�"B�������^���r�������$<�񕈮�3^8�8�>�jD-,�1}Wo��q���J~l���s��6��&������ჽ�e�ĳavx`r�WS��2�0��a\�'��@����RF�WF�]�>��n���tf�{�d�!ﳛ��5)q��%����~i���Ug�,<�EV:�|L�S*��)�>�aGK,)0�ϓMtD���l�9]�no/���e�&�,�r���Z��!o߷9�C2�K��۶�h3[���.�S�������o1a��q�R$7'^�ݙ��i���S2��5mg>���޺@ϋb�i��FF����glԠW����O�ʹ1��Xq�"H��vW�X�I,7�T��x�-G�y���@0�2�|�_���~�l>[{��ad|r�f8"�xS[Z��q�tt�Dz���>(����%�y�$m:>�o�)%j�S#c�(J�#�&M�ʆ�,WZ���(2���8�
�/~�__�Oed@��59:UдTa�k
�7hȍ?O��~F�$����gE��>�fO��wSU9�?:rZqC��-����B��u�֓��K�R��+�և_!-o��I")�~d����۹:3o��	�	��i�{�&�*�Ǳ,ձ�~�;
��~)v7���˟��9}l��R/:OA���_T1԰S��`ׄ�s�R��hHH=C'dsz0x|������u����#��������P�at���*��Ͱ�׷�HԗA�4�7Sd�.	�r�����Cg��B�&��
��Q�V�ÁC�شtyX@蛇n�1�F�#2��2n:d��Е#M�rP/�#�z�9�6)�8jr�|śL�Ȱ�S��EBq�_��3O=;*�2���սt0�Ț�&�ጦ�a�\�}�$p�e�c	���K�u`��!��x!\��&� &Dc�_էd:I��N[����ùY:�,!_tY0��,�?wQS�������,K�Q1u�#;3�`��Al��dG�:{clߏI�6�7�T=�-8�Lh���5�N׭�!lM�n��u햡���r����Mѽ����<�[;b�@�'+��`*W�r��@��$�)�H�Cc�,mU�|�[����eƖ�}�c���~G���^�JCN@�'�&lAS�C@,1��ju�	ό?��Н��ޔ�3���Z���?xA�����a�JCc]߲���y��f�<g��	��W�C�1���`]e���#����.!����c�N�z'�F�??+�bĝ� ��ݦ��J�zJJ{� ���`��ѺxM��T�0���x}�EPX�\�(��̆�qZ��is��"�y6��]id��q]�O����q�0��u�|��U 犿�u��5u ��Py���{�e�Yܰ�j���	A?:���>��U��'�Gϝz�QE�yI:f,���a�BT�O!�,�_��3�~�ui_@�lG'k�-��� �tq�ܛ�#��D�ӣl���M�M�!���1������IeY�Գk�$oY2�OuEK&��X��<I�Sj��NCH07���5#��E���Ȑ�5���g�x��t�-M ����hwz�����G�q��Wd����k��H�uy>�|���df�`��i�n�u�	�fA�C��3�o�)��z���^\�H�����J��08X��K0���an��Z��Y� $�l�����a^U`�l���>�:y=�����.��+J��R�Ðݕ��&�q!wy��V��!���Y]V+�G
4�t��	��i
�H3�P��dMdM��%!�$X�Ojs��"�w�_�Q[�.A��w�$�[Bu�����Q��3�M�';倳3\��W��v���� ϝ<�4R�Yf��Jx�y���H����z��-�m���Y�U,�2*/��17J�)W-�h�oG$M	/����a�{�� �ף��̥��o"^��m3��P�|�}���n�1���;7|��n��B>��~�W�2���G(�y��D���ۅ�]���҇�@���<�vu`b����3��/���7,c.h�ه8n�D��1���tq��ї�C�������Xm�͖2"?�Xw��LQXpP��o��-�>�x��"R�x�-pC�y��B�fxXK�>EGYd8��"壴�~W����*�"��:��NYdf#��F���>�9��<`Nnw�y�=�g `��u������H����XB��4��C�w��K�dd��M킜���U�M��YG%Ivhi�;�!����� �#�+�h�5��X �з�&��
��x؛HI!�|��r/~���0�?)��t�&�d�����f�]��k �<y=�~�}m)��A�0f�/�+_�-$�TU����6���>��A�i1&�)WBϢ}����L�ִ�&3dP|�N|�� ԫ���1,ϝ]R���ޥ�`�DA啂`A�D�\Âa9Лh�,��<O���(�s�Þ��.#˓�#��"�[��G�(��8su��������`&Td��'L+���'[oB��)yեJ�%$q}��жB?���6D�H�T�*�?�`$�X�C����5Ԯ��^�������i0�����K��hRA^d�#����N���ĎA*!�.5�ōX�I��5޷/�XB�}z�ӊAu�����@���X�)��l����	���]�nխ�=&�	V�E1�e�/��ΠJ)f�	�K��[�d����� ��fY����F�.EM��¢�h�`��kF;� Χ���Kef��d`&,0N�-��n[��
��'诮��1U�u����_�U 8!�o	��tI�M����. OX�P���lX�?�ז�2ǤQF�-���@�6n�V���It�e�`�e���gϊ'b�,�R���z�U9�i�6�8�{;��*'o�+G����M�����5�P�p�G&�J����m��	�?�쾽NF������f:fH���T{�Z��-Vix���v���|����Np��p
��0�����*k��'-���l��c����xL���_�,�q��"B�#�	�m�g��X�ߍ��$��2]]Cl�[j��G9����/Yh��v��<QH��J�L��H+��P_mO�z�F��d�W�u.I	�$���Z{��J�.95�1�yP	h͏
�;��*]`j�[��ۗ8��:`g����\��PW��2d��������Ds �v����7����7�r����Ӽ��^�(��K~M���P$�O��Q���5Q�$�˫s�uH�M��
8Ƹ�&��g����Bl�A"����ۚ�H��ibإ�٢����rc_��jt�*N����|�NIQ�������M@�9L_n��X����7��:15W����ƍ"�~�a5�7�X:v;�\%����h�1O�H7���Ĕ����N�����{����6��s��qx�����՝�WRw+������N��%D�Y�(p��ٰ���B������"oN1��W2�TR BH:�6)����;M��^�cٜ.o�c���G��D�Mʪ��=�ae�0�p����x7�(0��8'�j��7�,C���Yy�E"�u�c)@%�P�M�D�_}�U�9l-�Y�S_�a���nIB�w��=2�d�<|E��/*�``��M֓\��w���Ϲ9e�6��S7ɞ��Ǜ�+vS���F=n)y�TSƵ7�ܢcC78�Ҫp��w�)"E�[|[�2�,�dP�V�p��iO\K�t����)ـ,�Y���B�����9cӎ��0��p��6(���!� +�]g!� Zx�+NcК�'�����Q���мy��wO�jj��!�ӡ	�c�$�v�yx��	�qe��ҟ?���`�
������3o>JZ�[�wP������8��DrJP����̆�
_�L8mD�Ns�E���=<I�*�!M�^.üh;pT�7}UA ����
��u���^�,��¹S�s�DH2p�D}�����\g=��7��Y�.�7 �[L??�/�/����P��9�;�*��~x|��ZY0�	�)�A�L�� �Bv^�F�T9/?��bf��a�Y^A8�~)V�idʘ]�+A[pw�⟴BGf�-W�]5;y�h�*|[�����t q =g�ڃZz=��6.��^�;j΍�T�ÄȎ�><����)le��<s��J��m�^�ʢ=Ԫr^�.��B�w¨-Χ �NhɌ	R���=(�� ���qV�
�zo
U�A�^bV+`�T��z0�� X�j�=�V�G&OG��6�ЀR�z���)��+:-۔�ʉ���m"�E��m
�-+6S1�W���1����C�����xz%.�X�W�iZ<��� �2�ݥ�+��b�q�(���c.T��Ch��8%����Oz�clP"8���d*��=���4��}.��2t�<K�C��Z�v��<GD��y-�R-K��6��e�=�R�>p�����>h������JU�8�GPEət1���z�E������A%�w'�2�۾V�����<�4p���� M��������)3��)[�~.�V���V�a���OIؚ�Se���i�GA�9�'�@��c�0�>>�(��lAU��
�إ��8�z��tN�@�=V��}l�����74����;>�f�g��d�n<1�ՙ����GS���H�Ê�md����6�H,�����`y�ݒo�7{ <C�_���!��KI9� �GX�_{�_3�� �ox9l"�q+o|P����u�b��f�Z�zP�t���FK������0�6Q���8E��tϜ��������߼1=2���m��a�>PU�1�l����u�C��u�df$�����q:�Y-�D�F������3g\T��)~_I��P��)AU�����n˄���ų���mt�a<~��'u����';E��k� C���b�!� hڤ?nKT0F1C�5-��=$+��*����7��)r�Ԑ*��cZSă�tɒH��N,�b�Q����tr��kŻ�(�d4��rѥ7����<�X���&p#&�xZ�.��r(��$�ɢ-C)W����@rW����!B2X�2��D�C������]���0�����P�R����g�U,�P��a�80ߢ�6@�n����0�հ�G���ԘP�)k�kE ���蟰�L�k�ă��qj_�U3������&ұ�y�=��S�BgN>�(�nW��Ü��RfFq,���?=~�����F�~��t��q����R�3����\��w}�:�����<KB�|%���8Eh ���T+ s���vS��:Wr���K-O7xߚ�'�.N+ʉvW;�Ζ;a8��װ�˦�-Gn���z#�L�V�0K����1��-�-nEw_�=�eS��D�[U62�Ɋ�g��8�N(��G/>pw=[�p!ڒ4�I�c��lC`Q���ſg����0��H�M��c�\!Kj����3߾��U�[�'�y�9�F�fz�pP��H�_�4^�+�t����ݙ��8���M��}[S>5��ˈRh���tw2��چ�a�u�}�g�����>l3�b�j�GJ��2��	a�q��G�����D���c�i�%�,�h�@&�P����%\X�E�/�WC!\�S�����3��3f�i�uVN��{����ɘ
� ����ㆹs2�e��)
 aĮ.Z�^(j��7?I�( �E_,b�7Ri|�>!h4;>� T�{�jtJ'Z)rK}}���c��U_4�O��-V�!U��e
��N���{2Ìhʹ=��,��񶼮Q�	is.(�U�4P��vl�8��l%}����2p���ܖjreͽ��FYQ�Exv7#�D[U�~恷��~��R�CQchF]x��	i�E�)1@WL��&�d�l�Ԍ$�h�a@j�e�ˮ6�Y�ٶ_R�D������I���Pf�'�ݍg	��+���s��Z�F�����>�b.pdR�V��I.��J���l�+��᳄�`���=�E-vR�P�6���i��B�l�e��1��l�hC�C&��ߪO������߃ �_J ϊ\*xtyq�g�,Tj�0�G�@�ԇCGϧ=M��b2��J�{��VK��R�)��C��nDVd��	�QVb|����׬��&��pb�D�:A(��TkO�4*��5 �rr8K����.|��ҷ��F��%�!X�ֻL��m��w���l{y-aL��&�N�v�;j��Ն��0#q,��l[���RU�v� ��s��e�e�Ժ����m���8���yd3�)��&FԶ��Ԋ�jЪ��Z�O�2���,��,CW�(P��p�*e�&���u��R���f��s����HP�0���;�}�1����IY�����f(���O�-zU�s�L��<��PW����a.���"!�KQ��	�����$'�������RR���*��JnW+)�[M �>'��T[l൪Z�Ύ{H�ǬK�j��}�;q��@�@}3�o�:k�Z���l�'�o��)�r�3-��5�|��i��'8��C�����Y�5`�Oi�������5�/y/��
�bKz�^�u�΀����Bl쪇�;d��?�<��S���Z`�ߡ{�]s����s�Y���i��0\�C������˶�������2p��FI�3)K[-A`�>S(]EjX���J��КO#�C�W��$a�w����`(��>��ub� ��5v(�$��!�F0�|�v����N���y[ܘi�Q.	�-�[���R����Ή�%�Q���Mt�O��I��:ߊ���$��mKrJ�HD��㤁+���7Eʹ2g},�eǪy�	D%F�"���u#p ���J���Qk�ڮ�d ��!��O�D���	�Sh�k8�U�\�N��	�pd���� ��e��I'
Ȱ���$�^jɕ�h1�w;�5Q�4����.���m�n:;���'^qaN$#���к(� ��>b�thwqۮ&��c�����fr��4��!>->�)�$\�R�B�К��s�
Tw�����p�qaH�;��@�A�4����F�ݿc���\e�9x	執y���F%����e_鴶�XB��3=ͷqEQ�PF�V�_7H~�ì�&V�AX��G��'�b����PR)4�B.�Y�l�h>7h��AO�]���p�6����!:�p�O3f4І(F*C�=��v��Csni���N5�U!I�]]�2�����;�\v�+51����I�h���8V[�ׄP�0���o�*�۟�´鏽o�I�'�
�9�9�8��	��vyc�.B��$�#��Zӵ�P�-cm�ᮞ�W�v��2p�>��X�5�v9珚u�}X��LM�V�ӓغ�\VE��D�4rP�<��*=ȡ��>GϝGo�y���JD��*"5џ�5X/4G��{n��C��K�$",Ѯ�Cݎ�'���/ݚ(��	�\����tyǲ��͸�����LǸ<u������ĭf%YK�����]�!��3ϫ1>��l���$���S*6*h�M�y�q�H<�Q�:HQ����;�?����&
pd'y#�[����`?�|�����α�Dt��K� HXc�F�c�x'�$�Cv=�z�	6��. >%5N��إY$,����J�?p}�6m�W6�o/��i�v9B�U
����t���GR��r-uV�G,aS*ע�nuMH�r�F
��p�ڶbV �K���"�_I>� <A!�{-Cg���pw����j�<=t�/�̕S�P�
�����x����vV&�����n�F�����l�Vu]Yz�ǻ�� 3�9sp� �{[�y�~+��/}p����=h������tH]��򞍃G�C��zmf�^�o���j3��̋t;u�ug�m˺|}_�ӈ`!��L�a������g�l{���@�PȠ�0� '2���v�"��߅-m7 5R�T�=zr��;�҇�'�wں����K�Q���saw����x��r�-�"4���;A�]6�\��Ŧ`�ez.����Ȇ��x&�'�����NaSP(�	����r�$�-Y)֛�sV]��+��^R������[�e���;�=?R������?5+�	hy^��O�]�mo�j���^��<Hd��Å�0�&�_��9��D���,��۬��ܸ����J��>Ӄ,� �X�u�����R��J��d�1��� X1�t���֮��IO������Ga������E���NIu�^�����0]�CĹ��I��a��쏽u�f�k˻��_5hhg���C�hf�R����;�D��è1%:��vga3�/� S�TE]��� &��9��Y��gev�˳�8NZ0���7�*z*�
�N���%<:~t�*c��Q]�6�
��&��.����08yw��tg��^5m���l�&q�ɸ��<��]�I��
fu?Di&)��P��0-b�@��*d������U��'�ؾ������W�^����,XY��;��v'�~f&��{��l0P]�DPU��p��K�:pK�^@(�aQ�&	N�h���]�0�tգz��đ�N������&t~��q�[�·�18�s�XyPu�����:7t ���+�FE�EW7��˅��nn��z'-�Mm�y���t�����b�?oC��T �Ԍ#�*�����n����M2U^��z�_���΍���z��C4,SM�ͭ���j�k��](f@r���#���%��}~uV/��
y�rȕ�Ka���c���n������s�n��c��hƝӼ%�K��ۀ�-��W_$a����4�Ak?����I���yZ/����<�Q�v�,�F��1��+���bѝ���k�0�;�%��W�\��.�Q�O1�]tE����:�����Z��h�����6��p�%k�L'=(�)`�Y�`ColW�9de�``�t�5�q��~
�⃇ı��^��ğ&DvOb�`߼��V�IqmIՇ�)�;�"����ُ��=Y~�\:r������y�W�
Y6D� <���JWj��C!�C�G�D�3.��no�*�N$����9��N�c��j^��<nERn���!w˟ŁB�<uO��L�c��̥	 �I�`�9�>ׄ�E�t�i �%��B��	BafAKj������U�
�|�f��񡋳���[�އ�3�p�P�&"ב���خy�p��KH!ht|���l���C��K7�+$kz!-_��=��i��2��Gl���<_z+_����>��sѥI���g�'�C�t����V�$�����j�Ss�B*��@
�Q�t<iu�ǻ�"-哄1#������w��:D7M���(������k��L�ai6݉�����jҬ{��=�8�����Z�]1��T�,�z�T2E^����ڹ(@��oE˿��9k�JUaEY7���w^/�ޥ��Ȫ�y�2-ç�i��S��B��F�o8-�j������ȓ�Q�^��B�y�m5��������[X�� ��$��'�/p9�zޭ#��b^�u`���q�"ck5�2�Z4�h�oN��z���y2�+�p��^a���L�%�r&���o5�(=���DGݺ{6�:0$���iz(���#�/e��G��d���QFg�	*)����7ބ2!���f���Lʜ�^Q�(w��`��H�ȳ`��rsҿ5�mG�<�i�\��#?D�	��z��E�!=q�3l|�=�)�2�j@9��"�a�)��^�0������=�/��k�J�k�`���2�oFa	�V��I5z�b��֌���;脓ڱ��
=�w����Q *\:lª��x(�eG��{�̒h{�e����8��e6�I�y��
�M=T/>���+�=�OMsM�<'i"`b��Tλq2�Us�|�Ѩ���)��C�����^����T�mv����(X���O[����O O���نuV
��[��<��$�eF�Ԑ�1�I�0-I��U�3A�c;/�>?��9�����'�#�5P�W���MX<7[d~
5kW�A�-�Ku�U�P�}% �{sQ;P�)�lh@r|s�J�qCǪD��y�UV_��ra�ݶ��F�"�Ub�4\��*�XMq2�Q`'�ka��`1���k���)�4r��\M������7ž���Y�;���u }��z���y���%� a�F���̦ȃ�	Ro�R7g'%v��N:�����N5�W�x��z�X1L"�"�N`�C,�">�v�U����y��9���T�,,P��L�*�$އ�~v��B+����M������=D��bxm"�Ƴ�����DZ2��/W��i_=����q��:�*����������r�Y���'gT�)���鶅�kP�p`7����-��M]��(R17�,����.���v�O)d烏J����;m3/�|��.�2�,n�T�g]o�;����'������-���y�s��M\<I�z�W۸]��{�`2�M\�.zVg�AوƄ�� ���˜�����f��IC���j���/X�ŵ��fMKP���ؚ�n����W��=Me{��{b���Hi���[�q چ�Vz�Z�N�R�5�x�ER�~�:��m�R+�N��j&�����	�O�H�g��t`k��@�2HB������q �A�����Z����"�&0;�"�h����7�|�)���_��{(U�_�jKOP-&5it���GJ(�$�|�����ԛ���t]����������>�h��JT�;�G4F�K��E��6*�:���SAr|�N�M�$��w=���n�>�b�+�rL-�|&�`�q��U��gG���\	���K}�=6
�s\�ˎ@�� uwXL�rWt}�t������(t�s?]vY&E�T��ˑ���S�h4\��Tȅ���x-����
��揇w?�]q��*RZ`��_��>"�K8a/N'Z��ey���)���˔�� J��_�.�o����)�MwC�!Ϡ}�^iY*�

�c�Q^��J��3^��\��z�!�4G�����W�C*GRo��{�(��&O�6G"+u���c�'�	��K��\�u��p�`�NH�]�Q&��x�#��/�Z��е�ǒ����Y�M6�W�R|��~�2�=f�?�����V��:�۔r�����<%z�ƣP�QfZ�F���y�'|��"��x��::�������>I���=Cn��^��m���a@��'�=��o��qd�����%�����ֽ�zmJ���=��AM������q��<#�4��z)��q���zb6\\�%,e��Ӿ�j�<����ޥK�w�V$VL�_c%�j�ܤ�x	
Y�="� ��6iO���]w��}�T�����)@���8[����Kx���>C�W��Ƣ��>.��Ov!��X��L���l����۽ �0^8{ ��,I�v�GZ��(j��so�Q�e>[�/��-�K$����,'@M���%KB8�~EE�T-���C�|�1^�Kf����o*�9�3�� `�����+�1�!���lj�`���p�L�;�e��xhA-zA�W�/T�%�zh,�R[�_}��*Tн,e;I�K�p Q��'�-�F9HXhZ1�u���ݛ\7A�	��7L��a���y�	H_m?�Nj����1��#��#'Q��*�(=3�&=����g$p�I��b�^��@����K�)</�I\��ӗ"�غ�+�:���8��E��|^L6*�PF\���m)�U\�J�|�
�]�{ٔ^�P��� �yi����2��HMJ�>��dP��#@zI�g�D���kF*��Hq�ug4u�z�-�q{��8��ѩ��q�
�Y�=W޷���bЊ�k�1'Hn�����テ���D�ժ(��XϜ�N��R-��r����c�}Y��ii��L-�*��DGb
��Un�˓`��ៈ�@`U�� ���E=R�o�|�*`��[�'a%L���e��^P�SW��Y�ʆC�rK)�&�X�P+S�kg�f�г�qe"w��������YJ�F�j:��'�9�,C���%�a��J�o����6q-�T`>�L���O��0����Ca3!�L �_�}��>k� �@�O��'�f���bt$l ��D	���tv1C�$�O|i%�l�[�F�Z��z[z�;I�r���̯�)myʫ*���L&��dU,�GUF̧םS	v�f���úVB
 ���*	c����ꆮ�-��>���(F�ҁ����'ާ�Y\ljg��f���c$�j�u0�d�nJ\�$��)��`l�	�C lj�cɇ�c}�,8Q�ډ�}��&�ˆ�h݃�RA�G�r{���D�xNf�����7�٤9���G�%���ڮB��I�FC�b�zq�2&#R���<A��AI���R3�h�f+Ϛq�؀���U��e�Buu�Ϯ�
�V�Ma��Й"�����'h&�j��dR�`�C(Vs��v7���p��e�^��d���c��$�]5m��/[�5r�3�ʽ������!���nOH��fɫ�.6�c�u�b7�|�H�9����pg$�����#��2����Z��э�d���p�lWK�נ�濓s���z�)ۆ�m�����/X$�-U���n�Q��2up�3\@H�s���V��.O}�=����Z,�5􆃑���0��wa����S�7�;vbk�Yg	��=Y0-���^d"�Ī�
%���x���t�_ �t����!�es���<��52b7�C��ʩH���2���<��f�I�'0�Ut?v�����v�n�V�`u���#�Wq��p�f��	���F�Y ��������E�E��hj4��xz�����&�#��ċ=l���g(<䡰�O�����E�ݛ��R:J!�7�(��c��r{J/B�b�P��MmS
oLL�`$_M�A%�{��m�a�5 \��ZoG�9>b��d�3��ø]	L�i*�M��M�����7.)!�ĳ�0����t�4{�w��<��p�T�j ��wa:5r�1H�IT lQ�Kp\q��Ng�|�h�JU�ރ�]XYx��I�r���֚�:ڽc�$B8ܮӃ�����
�x�lF��9H��(D���l씆?|0�I*�e��`K�Ei��i_�r��1�Z9��0�g.����f�y�_�s9�� �k�kM�G��y�#Kq ̰��k&2� ��j��DO֋���"`�J�r9	��q�04p,�m����0#�G7 }8�b��v�t�3,i�.I�K�s�����dU���u��xd�1����
v�mR�[ɸ8�����+�IeXz�4�Ј*�K�
�tC�Y��ƃ7ܐ'�H�HHt�U��<�OB�tG#N�.�
PX�k�n��m]��耄�,�\K�g~��$�?�~��0y��?Ƶ���T�6��!3�����h-��T&q��2�3� h�������Z�	��`1jY��+,����%$�+������z���ne�A��~I~�U���e���'���#������&>������ľY�*C`4�b:�E�=ӶN��nW���>��*I �)S���2}�$t��l枨}O��@��+�K6cY�R�L�񶣊$:���96�y��P$E�B[#s�T8O�8�͈р�,͆U$C�R�(-?*h-����VK���[�U ��"T�|��2x_;�U�x����T��_�0�כg��ȏdĊ�#�N��u���ŏ�>�z�$=�x]A7\h.��w*��n�9<�'�/sj5v4qn�"|�vI�,_k����M"��%cC��B�x��U��ao�?y����3r�ː��|��q���k_鿍�k.ZҠ4`���S,.tm>����ɾ�-m� G��n�b�8i[;��[�d��O��������C].���+�%Y�)�D���r�����Z�dv�p�Ϋ*��A&�F��@X��aή�
� ��H2��#�vv�_c�4�z�7�+�a���,O��
gR��y�a�P���]]�)�*���%���򗫐b�r|�(|��)+!��w�L���}x*ݾ���K�pO��<�rȝ�ja~H+����됤J�-�~����e�4��$����E���Ɗe�_O�]eLeCㆸb(i���+�(���f5v���*m��"��b��<]��Q�{��zH���(�����+��uS�h��m1�!�&���L��-hv�~+Q�f�������ߓڛ
��	���^�T��0��ZDj
X"��N���S$Q��&DB\�a
5���At���A���Wc!D7�ʝفkxy6*k= �q0*Y�Ԭ�Lg�{�d�Hԇk�(@ )Ã`�:.�c�� q���K�ts�x��r���c�E�^��<�̤jE*]��{W��hO=�������,�'x U~��0��o����L��jYp�Dp�V/L0�3f�үY�,9?�(��+�߆�!�u$9�A�-�}�=�΍M�ߗ�b<ƽ�dD���p:�ax�2��/�ӼE���P�N�ge���NO���Za<O�r�Пpq��Z��;wW%��b� �ߥ�y��9Z�I��v�W�&he�}�'6ɫ��z�lQ}��m�{+G��� E��@�AW��&:UX9u�����U�sp؛�Z�Q$���S�{ӽ[�5Ӽ�r/�Q7�_���#��T��ӝ�T7�gY16ʐU3�f�6�rE�B����h#��d��U�}[�Hj�ǁ��x�����Ξ���]#YDmm�`�w����\��HP}�8K�;.�ݛRk�P���;:�l�@��k?�)s��B����`n�^��xttTxƉ�`¢ �z,%���{�oPhi�ceɠ�`z1��NyMFbfo�4b��k2m�C�r��p6k�i��
	�¢/J(�_��������i\��o
�]\���40H���Q��N5�O#��S�t-���A�|h��H}�^L,z��f�bI9ɗ*
�va�9����(�ƉFh]�Tl�:ȍ�~ѷ�)@��"�x l{@d��[u�E�@v�4���	����ɢ�U�&�KvycR��	H����{k�l
�D��'(D�.��&�5���,�s;�M7{[��߂ڙZ�����'�;1d��)L��0���-WY#�9��7V��\H�~��!��J�2��q�
��`JZ��r�-p-ՎMi�#�U꩷�Up]���!�('�=U�����y����b����l}�NK���(�B�0K>ERN��]��P��Z�*���´�r�g�#�\���ZZnx���q��J�'_
)�-�N=�ϭ��4L��c���`>?�$LB��u�L��-�-�K��9`N/Wa��Ag)ߞ�fh�B�n���}F��\.R�&�q�H�����^B@6�,�Y�QKy;'�S��8` `<�ǲB��fS�R�$C�k�%s�Yh�c��;�l�<_��j�]>�N;>��A ���c泬�{(vP{��ޫ��,��*���	��H���D���S�8�^=yc��oz�!V��YMk�?����d�M�I������8d� ��`��k
qrF�6q-�d0�d,��bS�Cb���BU_���,7l��;c��/�d7z�H�W�.�(3�q�p�W� sD��d����*��L���;�����=Z���)����,���=[\Xp��_�6l�(��� gڣ�`)��g���6$�k�ࠚ��=>+���Ʌa3����x���˝�P��uD�錹�����k�d�F�˨� G=~�R|�"f�O���j�j��y5���-Ww;������V}��T=�	`ڷ&ҁH���9�茉a��0�/%�ywhm���M(�$�{s�E v4�yJ�ӓn$�f���N�M�>PLd�I�C�na'��Bo��7��T"�e�pOH��<��Q_	:0�ְ��=�s�},3�H�?�6?�'���@�.�o�Ơ�-:Oi&�6�\*��H��S<��
!9���~���A!Q�:��{��2,8�D���=�
��H�4s6t�t��R�7�$.*�N`�r�
፩�u.�������:�5�E�n�.�ꁇ W�D�MϢ	�w��p7޹w��Y���*˿<łI mc��l��|�*��/�W�}7D���ߜ��6/:���	�ty�}Rer���Wp�0h���� �q�(��ԥ<sMD��|��dURZ)��t�AB�՘4#�F����������kgy�o��"к�����v���Z4�"�(�\��'U�= "�.Lϒ]g��M�~x<x$�F[�:79|Ϩ=y���4��-�T.mɉS�5���H��U��]4��a�b_����]c�#���W4l����]�A'R�q�;�-:t��1p΋f�G�)f8ԣ����n�@*�^��h�I��V��G#�h GL���ܚ�B�������fu�p+� ��;U{�w��zf�!L8F��%����ѕ��q���r�nZ�4���z��ñ���(��I�g]@�	���1X��]�_���$�������>O��C;�sR[i�3s?
�y,h�pY���_ �����/"�O�0i�m�ŧ_�`1��b9fḸ��U�C��e��W��C�	^����]���>\4�ސYײ���{�o��gm^6o!Ȥ8�'5��;�:��xأS�p����3>PX�q�~{�3��w���6�W��K�����.z����8<ԧ<��{y���l�⻵>F�)�Pwk���U�h	QJZr��S����B�[�{O𠅯�q�l����Q�/����4������~�&��Z׹P��]a�-"+���7{F��z�|;��x#��[E$���;��ϝ�?��7�1XW[FͰ���
S6�b��詬��d�-����+:���B�1����j���&�$/�,�&y��\��l߻�v̠���ݴ	��ֳh}RId�Y�����P�L�R�s)}�^r����8�v�������)܂2 >�W����&�jw}:nk3����|����~l	����{�m��"�T��,��q�����ஃ� �J�����'|C,���{<8�4�W&��Q�`[�K�`iwRC �; �5JR5G�
��[����D�O�@	&Xl�m6uk�Ī;�j;����*9�+�#-��AAnP�dQ��T.�k��Mn*]f�ν�1L�ߋ��[\����g|��df=�+��,�n>���y�����Pe�:*���1BVD��LJ}���Ct~9��NG�H_un�x�L�
�Z�~��ĩdG�+�=~6�G_]��,M򎂠�e�I�Ab 3�J$�[W����ˤ�y�]H�l�{�7�l�8�@�@!����Z W�����c����5�O��1`3S��^�� qkQ�Y��@�iڬ�֣6JG���pӡ�����n{�G�*����sD�kF��^'��V.@��
|@EίLh���B����ѿ1ei�1�B��J�����i���9�� .&�׵N\o��[[��Jo�^S�Jz]^�%kY���_ߵ��TB3��Su�nCEڹ�H�g�6�Þ�}�{��H2��H+�H���h���-�z���|�5%�I�b(�#h�8�`��H�ַL��5l�L����h�j^�f)�dAyN���ы
�C�(��E\쏤&�wD5��L�zfE+mE�w�צ�CD�%��rO�`���l����p#]s�)��6Q�ͼ�����̛o��,���w'	�P��O� �H��mEĐ��-gf�+�I����(踺���wqʇ�����H�хލ���u7�{��nl�?| �q0����=6ߑQ:��9���#"�%Y��W k&��qTJ�λ��)������=^����P.�5Ȍ^�bƹQ��op�ū�xx���6�8��S���
�&� ������By�����W�8�A�5ܮ�Yf�'�$}5���D��]��������� !���_iZ�d�/��yD���}���]�C$9�����j�K�E�\`<M�9r�"�j�੤�yn�[��.�ߣd��%�Y�7A�O����C���|:R��^9+r���4��i	��юU�B�ph��m�l�2�Ā�Ņ�߷^c��/�T����,�k
 �3�1!��g���-H�8aH�pN�Zq�\�m���]'���Z�l�ʉ�ޖ��@o*;᱖'�t)Bw�Պ�S޿�<�,f�sg���}�m�)Rjzef��� ~���фV��o ��M��~�Vq�ZF�ou�]u��Yft����]-/ޙ"���[�2`��+����$�XX���$��3����Q�U����u<���Pl[��X�7���}E�-t��[�Aw�P�}�'�.ZX��U_;[���	y�#�K�(bmڣdu� Yhz]�S�W��J5,����4	af'����;�[���~!�sC[����[���{̧�FB{5Y�]��3���p7\0���z�?��^�����ɐ���z3�ఙ����7���;0�гBnh�����Dj��D�ej�`W�I�s�,/7sR��+^��(������P���¼@y��]B����1��į	j�KM��I�b���l�Rb�Xz�#�2��3�����c�75�.eK��?�aCp�e]A�J6��4�ܪ5�C�m$�-�ͮ��a	f�\{2_<��h`���Q�m�$�P�� �� 
�1�	̰Q��d�:�	��؝rq���%�o�Ф�$XAX���"�5���n ��`H��W��߳�Ҟ����߃+��&����IQ��b5�B�Z"�פ�{�$�x7�t�`�1*���yN�Z��a)M۪�*ϲ��\�1�:�R�Y��L�r��U=4��e�RY�%���d$d�����;~���7|�GOom1#��i�<�V�ԉHi�2#ͤ��h�M���q'�ό*�8�B����4D����Q��
���4���6��$�mg1��e#�,�sW��Wq��ce �0y���/��i'>�f���1�)]5K�f:|s�8E"����k �\4�ͭ8���46�C��0B���۶'��u�!N�8S>w��2���
5���)�ձ�%+�z�f��`}���f%��s�z����U��MC��&Z��1EFdܶ?�������{V�jP��7���I�9�ܽ2�	oQLzj��tv)�U��T�~����V��pW�O���&
Rz��D��2�{��RK���p�B���U �:wf�d}[�K�I�J�x$7��mD��D`�߆T#<�k�.Wp=��&�>�f�'O�=��}'܇&�*��1aW?�C%�a)�D�z����g�?
�E�؋�+��P�ǆ��7�L�va�Fΐ��P24}��#���d������ٱ��[R-��QI�%w�0|�M/.�h�N�q6��	��B�"�%��ۆ<��5�iZ��2��pp#9�=��8��\K�L݉/�����pkB6��Hv�U(ߑ��_g�l�ƛ����/������:=:�6L���*���R��<9'��tL���b+�t1��@�4$Ā%G-!�E�<�E��mh-da���䴮�� ��J�h�~b ��l��Od�;5Z{�y�kk޿,Km��9W��h=��t{,GNaq�K��Oy���Ϡ�v���5����wH`LGZ|�JG^_����ވ��]�9�"��[�Ao�n�S|�'RԹA��1��W�n�g.':=J�8��'BվO��ۚR�Y�%�Rn�����T�5ށ���D&�Ϗ�OZǴ�G��̧h��
�\��U<�j)��&�K�������ti(6���|�3���*�!iW#�)�f��b�+�πЉfЍD"ir"���\T��R�'.#{A���	��kQ!��t�W]K�ꎇ`�����2���oK��V�J��.��F۱g|U�|S�j=˃��w��,:�<�^�C��½��|�r�Bǖ��,��#�\&5�xz�}SI8���E�;�l�ȟSJ5R�`Ҙ��lB�yT�y�ܡ��6z!d���+0��s�
K�'�-��Swwx+�@�D(�♇�o�\��>�`Z��i�e�V��(���<�1)�W�+�~'=Č�o=Aa �C�hj��X��V�/��I��Ӿ&�F0a(��q�j�����O�1�oV��l�*��0�<t������;�(�@�h��x7�Q�L��\75�:L37�j�;�������7m7�c!�4���2k�e��O�L	1]h%=���7]����:�����;x8�jsc�=�Ӱ���#C,p�gl�_��b�J�������Jِ*�;_I�y/�I�EFśFG�o&�ܡ��x�4k�m�Ԇ�G'�~�$Qx.��U��.3��}_�$�o�D�\���;��Q"3�����j*k�."��ՂeOj���`�\�obmA�F�/@�g�x��럸�Io���Y���7�`��E֎nW8� �Ϝ�p昳͑�������i�)�]�p��T��W~�3�2k����}\Ǵ���,<��:2�Ꟑx^����,<����dm^�<�BÁ3����x�TN�A�z(�+���z���|c�8N�2��CV�W�+P�a�Zд���8Xz��Xr��Օ�Fec�p�s�����u�Υ�ZȽ��~���:����[���
��ݤA g�k3K,���ZT*����'�y��a5���l�����jǜ�Ճ4l�1�ݮ�4�N=N�7��.�y��d\�Cw���<�['�)+�}	����@.l����p���l��Mt7hxf��Y�nkE��� b��#?!��F��W��?�e#@��8w���<O��Q�u1��#߃c����DP���m�']o~DXܧUi{y�K7����ۦn�:='�&���'V�l:�3eݻ&z��i��mO���Xk��8���Z �K�2c�]���L��Vk[�5gY�&f���"&�q	����L�F���ۿ�9؈� ��A<�K|�iMB�0~�{���M���� \���~��|�����->ES=�0,~P�%b�bq��&�p�ЂlHi*~R��8���V���t� �j؁��&�uHS�͔�n�N���$欱�2���l({Z:g#����ڵ�,�	Fv����<�#8��V����O�;�-~�͹C�Q�)�����Aa�^��j���L
�͵2!�Y�DRd��j��v�cv}Z{�N��b6�K�<�K����EN�g�����MQU�Dc ���>���of��-� ��R)$�a��O�u[1sK�X�S����vIY	G����UA��J%��:���{b(u�{qVA	؊���M�^��@�ϵ���J���>30a �~��̈V3�L_9��ߘ�ϗ�w	<��AG�����)�F�_W�kq_W}���RWW�ZZ+jl�
�~�M
#�܎��`�%+l
o���i����#E�O3��y+���)3Y�_�]`鐋���CFu+�l���[QS��{Gq�|�`~��&�*
u&a�~�O*}��ӂ�����հ4�B Ѳh��;y�:����M��p��뛊��e���A�����rN$[dJ81Kx�T�G8� ԇ>8�����!ǯJI�!n�Ƃo5uʧ^=� T�ga���t8����sK��=\�EO���?���9-D�����-rY|hW��;���obp�����~�02M���buZ8�|�Q���/����:��W����� 5�P���&�;��W$�ݜ���L [z��BX?hL5l[��ea������em�c�b��l�2�ŉ"?�����=2'�A���p�=6�d�*j\��U��울f�wRƊ	�|eP�Nw�J�0 nG�-��<��r	��Q��V�zѷRo�C5����k��d�8q2���������
��3X$�}��忡r�7`}Љ�jB�#8�#�L`@]��.{5��/F���9���I�Zq��"���5�s�C������J�E��-�K�>�≤��")4v�]�͙ݶ�`軇y��Ip�ĊD�ǫ�͒hH������C�&$� '���?��۾ ��4ض5�'����w.{t�+B��/yn.?�-	'�%0��k۟�����k���ح(���|��;�C�93�����������6��0fh��F	�}@�,_�7��&��Nb�fٗ�����-��s�7�O�i'�7�5�CT��	BU�Ȓ�l⥛�}|��&%�����$6�Ŋ�R����]�	�܎}-FQ[��\ʭ�6Z��y�����N`V�d�Pԛ�t�d�
�{�q���i�l�>��t��_dَ�jF<_��}��g�&1	�O)nz�'#/�FånV�/�#�l�~���G���\��������8Ѵ���H��2������E�i;�����	c쿤݆���@�b�;-j��q�zk�C���tc�I�c���{�����S~�{;���ߔf�'��mm�UcN�3�.��}Q�օ���#�>���� �z ���Ov�?��<����&^�rό���Ё�w1�z������.��P�	uD��B�0�֎��{��}���`���[�U^�djR�Y!�4~.$u\;,c�骀���=6���V�y{И�y���9�l�Ð�yuᾝ���k�9 iX�j*�� ���w�%�J�ԩ~��m!�̦�iE�5z%�u���d4��n!��KI�@nTi���f`SM��a2�iW�)�>X��1(�����'����l �L�z�W��~/�_��4������ӝN4w��'AS��r*ˮj�Se#�3�eP�W�k%`��~�I��%��¤���gMc��˒X���^Lx֞��@�s���ϡ�O�+P�,w�ì�*'䢀`X�_�jd�8�u5\A�0��Q� Z�l��	O[x{�r���\���I����;j*6�Ɔ��հ�+p�m^���Lg���f�A�fi�KnS2��4�Oy�+�w�s����I��/�eSIx@Z����j��V� ��ⅱ�ռ�QA�����M$�}N=eQ��ʫ�J�.8}�.��v8iY�p�xvR�:�1����r,Lct�/>=��I�W݂`�daD�+?�6aLi�a*�G���gG��e���{	>����C��犙47R�3�#T �F�@/`�ȯg �x��e��$e���)5z��콰����/F���J��1���^R��1n���t�b�r~J��3�o�ɻN*�:w�{ר����1UƗ4GOót�������Ά!�O����lsß���j[�{劷�Ϭ��ď�y�)/����^�8B��2�]��
{���kͯ{��?bx.1���a�?������NS�+k����'�U�};22����ǛP��#h��@ᐟ���Ўg��	 �"�����9�!�v�9�b�q�� �32�ħ�ɟ��L���g"�U���+��c�Y�2�s�tl�ܽ������T��^�(9�|�R�(�X�e�1���}V&��9H�b�a��n>PM����)���lN�q�����Փ�4OB�%�o�q�nOW]�-~1� =�G��1�^�g����/EP@R+�n���F�pV�������82��\ۑ�	aù�π��������ļqy����Fz������d�//9�,�?E1R �b��q��]
� p�]i�cZ~��2�[/�"�����Jx��e�z.F�	_��=俋�i�b3��y�w8�aF�B����?8_ ���O�q|�^�x�I�~�E|)H�~���Z-����B+9��:�m/@����#׬4�y���.X�i�L�a7��|�"H��8�k���ǶgC�H����ǪeC ����]]�v�Xه�u_��
"�δK����C��Z��v�o�y��:�{�\�_�~�ͣp�FX-jB�'�b��Rilo�+���UVi�?F��Ç:ƀ$��	^;��x�ܹ�F�rQ��D5�˷{�q�S�R(�Xe&��m��;��Q3������=�� m�b��w���~0
�nu�ɐ^�l	J1���D_�����K� e`�_��F�VNz���=��'�VC2�b�>�����!Q&l���I�;xN^��b�<2(kT-�!/m?���W�\�������h<�-�V� ��P8
K���y�60����$�]6����,)��ail<P�[����nR���D�ϣ�Yw��<S`�&t ����c�]z�"��-�$�b���wW3/�R}6��#zN�GE���5����� hN�=I?�B{g��N����}�x���H��Z�](�:���Uc{��s��,^Y�C��zr���:�m�a�������h��!��H"B�pF9U	�ӆ�m pl%!6�������������5�Gj�̽�n����q����6�L��K�u�S�M�
h'�h�U!$�l�j�/r��������e"�2�X���&��eݕ�
���(4N�d
�kJn����U)���VV���Gp�&q�>M`�R�HJ�\� iG��62�;��z~��Ќ�s}k|==2L.O���x��B�;����Gxm�WL+Z��ܙIA���V��a�mY,K܋s�Ӡe�� U��i��?�Nu���� 7���I�[*�һ]V)ZP#�ٛ���VL��n7�i�ڂ����ԓmэ���q���62������EE^s���({����������'�M��MX��	B�:+yCL5��[�f`�l����)��<�U�8`��6Q|	��侤�Ƃ�������!�n�� ����# ��d�G�.��I�.��^���+�Ŏ#z��j������]���A����=%z���[� O©�Z捾T�F4��0���,�U��_�?X��Rb���� O���x���H.��2�ش�ꥠ�{�C���6�8���4>U���u����m�g�0���~�@�i����O8� ��d�R�[����E#!��;��Er���ui���������+_2�C�G�23����	qJ��G2M�^A-P9}a�����`�^gthC(.#���0��&rQ&E��l�#�v]GB�����R@�M�U��������NE�i����)�O �\2�_"���:���&e5�˒�6k��u�.dű�U��^F\'bA,�� �X#�*�?e����Z�U>��-)8?ܧVu��S�����Tȯ�K��fVI�We��M]h�8���K��C
éX�$gص��Q.�������Nz��M2Qp�LEE��Ζ��ϩm�kT/=g�_�t�ޥ�J6ۧj� y�h�}Q{o��nz�O�+��������b�I~�\��1~R�Q�<�.�&h>:/��~H����o�������V$^��ß�O�`�.��H�������2���ru�s,��ab��ҹ/�)sj�/�Q;x���d�A"��w�}~�(��{WP���.5�_Z��Fp|��]q��%)���w�Bې�/��8��R_�{BM1+��<?�@�� E�'ͱȑ���)�R������s�Zt�wT�W�:�+؎� ÕpM�fO#�G��|M`����*������H.����V��ǩl��W��{gJS/u��!W�������ӵP�+��0���یS�#=R�+J�2�rDuD�A�m��Q���@I�ɅV��k%����������"��Qa��W��b��JF��B����(����'ی����TD�3��[8�0u�Ϩ)@�ߙ�q�c^�s��D�5���a��0��l�<���� f���66'�k�Rua�/ӭ��'� �|B�@7��/5>�������}<�[�0PeM�݃��Qp�>*��ؗ�2w�:�߃��-���r�Ҋm]�l������d_���ç�
�#����M�P59�\��fye8���v,�{o�K)Za̹.Ao���]�Ջ��;�ρ��>�M��������\�..8A�,H�{���/���K�s�@�`��I�C�d��-cOl��a�O��3��Lp�Y��k��Yb�6.�̇
�	E�!E�0��W���"�ѣ��mEZ��:�0+�A-��L��Zs��kz� �MT� Nh�܈��TU�p�5�\3mc!Q��53��vM�F�cr�%6��k���ez�l�q�/�l��f���#�����1ҭ�~ m�㯺�.!Q�E��P�A���X�mX��{�����	��|��6���.=�det�;g���
���cJM��*j�^3��A�7P4Գy�����<����ԑ^�v�� �a�.�"����ց�>��I�ٝ&���N��~lR��^�_Ի%�x�̞����Hq�S�lיִU�dZq맕��۾�\醥, ��>�� uW8[�q����g�v3I��,�-�R4�:�Џ����r�K�422�w�x��S��j�6_?�(R��F�I3�piҥ��1U ���b L'���cϑ�" �	� .�{�Y�A�l�6�\����Dc����j�3t0�24�&|1����J�Ң S|P� 7���d��%k���H�m:��Y���*�fmTF����ɱ5@SDlB��B��C���n"�wȦ�NkBt��Z��`g�s^4h��|<W�l��r����1�Pk��� ����T����W]�P�o[�yP�G�g��N�����T|amS�db'ݗ&m�r�/���8bK;�n+p�������9j�ȭh��(�2<�����Í�h�:g��\���%=���#2;o$Π����/A��$��|E<n�
�R��z9�,t��53��7<���@�����z՗�׬��;l�΢�+q�F�l_LoD�C��ke{��!#���d�2�s��:��3��(���h,�ep}.Y3Z�^����x\-��f��E�������M�q,DmD����E!m�n�m�(?��+G�E�
�䔶��+�t�Ӱ8��'��j�Π�jlށ�w��>��uNK�^��#㳯�W+K��(��U�͇8�=q&
�Tu詤���YF����"xzùk=e��=�Ж���w�����'�y����}��XUTYj����K��	pZ9r?pR��*�Cq��H=� d��.;��:��f�lT�# [(��g��n�:�Z���I�"��O�oL�����R{�>�7�׃q�Il���rpz�v$�7L�S
�
>d�
6�G� �QG���g¨z��7�M��^7��� ����**,F������09F��7�I��kf�v�$���ڷX`GǗ����j|�Y"�
j�H����5qyQw�+�;�Q�0"E�,���	\�X�3�p��r�1#��5Ӭ1g����0gN�Į���_����}�cB�;mZ��S��AeKe��"JB4�1|QI"獅��¢Ͼy�R$]i�5����nq�!���酞(r��i���$�������8U~�5< �
���nVo���Т̱���!��;�Wl��Տkb�t�� �g���&��\jD$U{����U�ņ�N>6H!0���r���vz�.,T��V��K�6�:��3�g6�̏)0����d��u*c��,ݧ>4���]_SxjXe�qr霭:��I�ȴg�|Xh�M��(w�&{�2IA-��]�TI#*�5�����w�~+�]�|"�N�k���4�*��!�ݦ���T��6:�����0��u;�r!��l}T�ެej�q�y�����ĳ�p�4�=��k�l��^����ٱKv�����@[�P�K��I��=ڸ`�d�����S�e�8��=�_�ٍc����WR�͠S҄�M"{%�nO%O(��V�j��RӒሆ�Խ)7#�T�u�LNڏ:�
�.�} ήM�"�y���(o�l#�%�#�\ĳ�I�hv��wS�&�q���<!��$�����Δ\�{����k�D���%��@v��E�����#��L+�;��	1ݫm̛�2������J:��:q;�#��S�C4e����޸�Qj��oXwT'@PMF�R���F�:|�l�m ��BNk5�M����͞�b#q��r�.i�_���`ыT/�c)q�8�f��
V�]/�N����V�t]K0�S����*�T�Y�5�����y�{`�E�[�o���{�D��-�A�کB���}�����2{o�`�J"g�?v�l�����3�	�|v�'0�5d�t�q���K�i���ǒu?-����˛���\koQ��j��ދ�*u���pr����>^��AZA�Uw�����	��u[L��zx'�Y���L�eG��Y��ʼ���Z��~���|v�Z���ir�����B�Vu�w-�5^#g�F����r�O��}8���j�Rlk� �'T��J���3[4~#�^�vE����w�(y�7�����ؽ\����7����Fz��i�%`B��������CXs����-^5�������y!�ړ������M�-A����O�rr����޳|�燐 K0��M�Y���Tw��q��
�0�2����X���<�M��pg�݄^1�S��M�ޕ��73�)D�[BN���W*>.���ɓ�
2�/�ľ�Z?�Dy�[���%�.y�~��w��(��;�q���gck.�^W����b�B�g��9���1�BT׸��N>�N�s���-���b��˓�y�q�|��k$���L�@_��%���{3���O�yNӜ�H��|���5Bњ����0iW�h���J�"%0c��?��W�Yh^�"��zП��w���^Y��:$*�q�?u���I=�v�&�=0<�4<���_^��Th����*�%	!��
3
[�S	〴]UvuE��{	���.�n��
�pg�c��Йuٽ�B���4�2��5��`
FJ`p���:	Ɣ�_5��v�)�#ޅ�b���M!I�U{"��� HT�0�ը�4�V����qCS��z�[�v��Z�3��*�U���*���ל��TOU�v,�y��r���o��������A��pH�ԯ�s�ٹKGNC�yg?L�ΤS�C�gA�H���b�0;#>U=%O����-�%.�H �1�<.�A&�Z�n�yJ�9ü[��0��4P��]IY���E"��_x�����I<.5x�b�F�0̚EYP޹������s}��կӭ�ƈ�z$��Ch/Ii���
"r�[����5�c �E0�b��iyi�{a1k�de!��� s�:\H�b�^T��y�ϒP84�Y�����L��2y�Gy~=�� i`��=��?�Zkϰ�53�0P�C�pM�����Qi1KFxJͦ�n�}^;rv��kJF&���h!p���-�TM8�h�����{o�\v�xrVb��
�՜��h�yF�+�J!�I�b\���⽐d7���"�8�f,�)��Ċ����|������Pѷ9MB8xj��L�
��)�j�)S���}�t����^
� �~LI���jx��(�Qr�Id3�Aa������ ��wN�ʲMX?6��Q���<�S���|RpZLJ-Fdw����]A�c��p9
c���"V���n�Q�w�H�I�GF���($���^qT�x7�"UdpB��� J����7�<���YR���Vy}�n���V(d�tq�x��2�������=��z�b[s��&�����a���z ${��6��GҎ�!��i�/�,ZɄ���'[�LP�/\� ���n��-p TB��6�M�k�0�c5����omέ�ɝxm�ģu���.�a��F���{��{��V�|{�%x�����p��%��7�&�ګcA�5~����q,��5��fp�vEIDM�jzx����wQ��1d��r��V���> ������"��I`�6�,;�3�u��$N���L
6����=�BxA�f-kJ[�g����JҵEHș-���S�t}T^�Cg�N��]/����cc�)=�q6OZW>	�{Q��TG�DQ������3Ɖ��o�*��M�NgV�9�;p�P��0��D 일Ș��p��"������l�g4&hȕz\�W}��な�G}�&]O�>%��,֫p��T'	��CX���#�@{���Uz�V��Bz��)@�YȧNkl�h\H$b�ދ
v܅FJ�p��BR�K�'`(��V/�M��K�萛�J�]�в"�P�Ӊ���4� �6!p�݃/_$�h��kg����:�nT<�^�$@�jo���1p�ŞC$�9��Lt��#h��}�gГ���Z���2���(	VkQ�\�hE	����P��b4�;�y�����楬��\�a��d�0G��Y��U`c�:R`��j��|7�l6�1���u��X�x�I�#����Y�H����-4��` �iX�{���xU#o]$.(����lVK��!d2lf�W3	���J��K����c34x8�r���bb-oGg����p�<NF�}���?lc���:��>�wT܏x�����q����զ�Q��B��p3qn\�9ۙ�leN9Λ�\3�ধ����"uE�6��"�Nݰh|^+yi��m�W.���<���X~�������A�L^�Q�Ϙ_������m�&'L������R�����ͅ�������y��	��aO�̰Z	aqP�����(�J��L),#���3$CM�~%�9o�S�C��.�yy���˂%��c\���{nw�닠����)h�/1n��o�n�����mX*���8 ���<H��nƅP���=z���;'/��K��|��v�h������ϴ����
8g�=��;�ʝ6()W���7�#�Y`����B��V�!k�
>�]�'�fX������3�Sصrh������L��w�C��J2��rV�z�4eBF�i����t�[��G�o|}�@����T�S���^i��$��j�3���NW�k~��[��Z;�� �ɷa�D��e����,>����ћD����p#��п��e��Ύ��ɫg� �E"Ǿp�a	L��`�kp(,�|8ˉ�c�,�v�o�{T�g8ح�����;߲;HZ,Q��@���N�q0�&��}ج��$�d"	��
��k�I�
����o#�x�ô\�K�/O�.QN�\rW�I&�������R���lH����r	:iM��!�g��/�^�x��P�ºyr"��uхr�=_+�!at圤]ޡM�����]ߙ3��_P
����
�$H�����4W9��,�Z��D7�D �u2�uw#|���`��1}v�����`�����x���~a�$�\�=f�Z&Eb|��[e5cԵ�76Q��3^�2D�h@�����_��/>	N8e��c	����5
��0���"�
�ڃ���j>S?t}tpuH�I������b�M3Es_��@)���C����{�wU���þcw�y�����̗@g%a����|S�z]�S��z�����L�xb�M��d��o�Q���3Ȧ�>��K��Oco����9}x�m�F)��c�_2-~���q�7j� �����Դ��}�:�L��aۦC�us՟4�v��eS�j�.%v?.��$PeN�s��s1C�՗?�n��	�.�T���t?nȋ�Q�un�Q���'`Fcmv6�4��'��U���4�
�8�#me�P�t��Nӟ5E��m�����[$��џ�!v�*J�-T�Uwf�}/�� E��V��-6q(���g���YK��E<���)���t׽���/[��\�{$�+�w�]��d�bnƯ��z�C�[�=���n���y���ݢ�)��W�2P�i�6�/\�T)�a�A��lq�~�Ř���j �M��I�_�IWH�=��{�.�j7�<ȯd,5��S������C�bYDW��:S�v�<<h�	T�`q�ec���ԑPg0��X����p�;��;���DB��	����xq[��d	y�u���Y�z���8�ܷ!xla�hh%��$�/P�)�/*=w�:�7�H:e�G���s*�9���V�H�&$9Lm�S�_�p��E;�r�/K��m)U�ߜ�P#�a�9g�ui?
І�vr���o�8p\��@��Q��'p("y�[,��(���s?�KCH����>`!�^<Q�*_���%5��$G�5��zm�-4�#Z�L��~��]�ҍ�SC�s��]�Y����R�F�*FH��3OU/�L2�X
��kwU+4�]�����,���[-p�"�7W�wI
��d���$x�$�,MT�_T�+&�w��} FK��\&I���KP\N��]j���`�1b�AH��I�ف�����<"�Y$vOa<P�i�H�i0�}w
��B�f�Nm(���xJwWP E�	�Gf�# 	�<�ԢR�[��s���@�ho�w����X�>�/ň��UEzTEh�ŜW�t�n
h�
jj��)V�l�?� -J��n���.��tTr̛xD' �bf�{�����c�Rw���˷����˔Z���힡@@����+.R#i����PKÙ4���*���J&�DM_�e�1��$eq�����Ns���~�o=��)�}��q�cG��2�7�,g�����*l��3� U��@�_Z�T���8ª�D\��k��+F�{�B�ٳ >����=�	��Oe��PghX�A1�fA��E�R��E�8�q2����~�&��x앢b]��[���T�[�߮^�XY1�] Ǿy�w�VB�GS�4�!�x��H�r;��A@"'�J�K��1�r3�XM���ZMknu�y�s������b7��V~0�[ۆ�kH����������g/�$�s�uM��%k�w|7ǷB	T�����j�Z
�˜�R$\�����{$��_���%��������"���z�)��xF�*���jdvD�j����ǎv���7mC>>>Ld�˺v��� f��<��.�6��|�o�a�Ϳb}�����+������+���ݨ�t\�Bf�	�N��f� *�����u\�z,֛>�ԅqPR�t��te���i��+&ݞ����w�x�xfBu��#���6<P��h�w/�	K�5Au��ҳ{�����k� �9�|������&M�B�L�b^R*�M_e����3(����1_:Q��6��"wW>��;��
X2����jn�AXP-�>��@����PԒjcBכ�h�&o��8���UW��a�V����x���/ą�b�6aK_�����=�7TX�"����F�
�^�E����j��#l(��d5����R��7����:�"�o^��l=��Q�+�~���GX��k���7ʱ�z���bv���J+�>�F���m��գw���tc��e9^PHM��G�`�
��aB�~mQ7��ׁj�E��J�J۪�I��62L?;>q�1}��"/�&QO�k�Y��Bh+C�	�	���FT;��xy�R�
[$�~YH��̛��>�k�����?��Clg5��(�Ejn��}t��?6��8r��%�e1�ϦKY��Gֳ��rAP��Z4<�������l��k����~Ap�	�q�+Sv�4��cg�o�9�gڊe��-flbs�b����x5Y�/�%�<0V&0cj&j���2R-HEM�ݱ�O;�F����/�qb{n��5�X얄���`�d����5SD.�:�����E�/6��O���'�����9@d�uӭ�+��·?����}>v�zr���8@���'��6I�֦M�͈zR� <w���\��@�Js�H�m&�y{&.#�y;�"H����} b�,�.S���A�݊�m;�
�������uR��1��|���z��	^�u�� ���l�Q[�w˄��ْʹ�`��)�$��pX���{���nj����W� �`�r��<6�:����J��{/s}\�D��������7<�?�ڹ�����)?,��N��+��L/7��:D������|t�]|��[V�d�����R#	��'�i���-9E�4�cκ]T��2������ìo�c�l�dI�C<���x�)O�Bo|���kr���r�i���v2��'�=ŝ���&�%���.�/�燪Aܬ�NBjY*��r�-[�W~{8��\PL��Kъ�H��TN�f� �SR��v�Wc��ԍW�|� ̟$E����>ۖ��� ��������S�ӫ3ؔ���,nF�`�d�k�6��7�	
�j�����P�<2"���]��((�3�$�hX�8���H~�����8Yg����f77 ���1(LV����\k����R8~�z�����_U���Q�����\z+,�|=U�JbkK3}�7�������>��b���.�Y���?�O��������L ��[�����4��c�u��^�\О��=/��6[����>_�������ﰪ�IFs�'�^7 խ����㤧��p�;� �3�N3SWF�z}g�j?�4+΃�lS��c�������#�-q-�J��>�>�6�%*� =���%��`IuC1^yL$G���+Oq�� �b�JS�z�#���V/�}���!�k'��6#ۯKA�
�酇L�6ط�2��9��:4��h�UXZ����qjQf�����޿������)����R���[
<�iQ7�!��H�����Ydwe�"���e�������}C;�\�?o1��e<h>~#�.�ؕ��v��4r�!@����;T�
�����R.9`KT���py
TN�8Ǧ5�:��ݔ�K�g��e'&�S���D5��y�^�����Q�5}��[�bM��]��������o��UB����+	`]��@F0�����]�H��R��Q�@�=� I�<M�+ݼ��� 56��%<�  �� �%2q3Jr5B�S~�Ha�?�bs���QG���Q�7��<�IԖy�"�;�]�*f�2i�F�:��V�i��A�ߗIxξ�W��5��yY���a�L��e��W����1t��R:���|�~ �d͂t(���oj�qùķ�D}�l��8Ae�����R�i���=������`)��L^r8�-�L��<�:t4Y���+���x��;�Nu�3����*�7�:J�+�R��!�y���6�ܿ#�ʺ|A=rO��t;mdP#�le����5��^-�Q�vXNy$ۙ�i7xw�P+��_o'��o���ʁ��=���F ��O�� ����B�p�S����Zvٖ���aZ<B*�7�d�x�є�`����R5*���.��E}�j7u��8�J��ⵣ�>�������)�N$���-i��lD,�_���JI�l������F�c�l�솽��r��p&�?!��LB(^d3=ha���2#&ї��[�an7��4�F��+5]�[��I���޹g��R䱸r+�,����[�����|�i遺+� ��X�q��fI�TVm��r�p_d8)
�>�G�b��n��9�2>�.5x�������K�������|D8�W�j�eǗ2_d�`��93DyG�J�~D���_'h��t���ڻ���Lߍ���K)�P��\A$cH�]o	{�N �/��ˆFG܈�-j_v��G��P���_�h�͗������$OR�.\�fK�������G)(���.|�������\??0��d�+m�b���C�x��Í�~ϝ:`��v��}5)l+�a�)�&Qȴ�[F��+!�A}������̲�SҺ7�\�QC�����M�B��B����_�,<���Vl�\F�=�Q�R����GE�׆��o�7���0��_{���𒵣d��-XX��ǯ)��ְ4�M�Lʰ���8��B[a;�xg�0���)"�4d�g	�aV���,Wj��������@4!L�륷2�.�M�Ϝ'�|�+�)�!=���;��A���,\�[[���:4�2��%�l� �MSE��<�Q��"����ɓ���d�d�*b�2
���e{T��j����L��Ջ��D�����l$�	�*-?���l�S����{?Ӽ��^�9���6m����C7׸����#z�������>��sY�������̱Z�$x��^dᖒ���ڱ!Ƃ+.��}�O>��_j�c�Sx\4S�>T4y��ݩ�P�=��&�W]v�u�a�u5�R��S��NLr�^�Cw-�@����a��ٹO��wN�z��j�{'�!���e�@���&"#o-a���~š�Q�0�킇���xH/ߟ����`��`=��8.۵"V���~�&�,��gE	�
Ҏ��tK�`��i����#��#��� �����w�P�h��I�vt>�q�n�-