��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%����:P�f%��mnn��Dm�n%N�w
�cM����_�WJ������Y�G%Ih��|���m]�)�v�v������ք�jc��⾝(�����Fh�.��m�6�iy'�m���)��V�����aGo�����Nh+g�lք���`�l2�؟˪��Jh�Յyok��!����8���)�� �CЇ��N�d�Cy�X�g�&�=A���cS7\�����s%@fC��j���G=���ܽ�P���������9���r삾Vi�tC�;�A�(Y:l����>���5ݐ���9��μ(�Q oG��8XY��RQ�튲L�rfpw����f�L�u�W�')C���Gڦ�z�	9��@�~s|��xs�;���
�3�lL�K)��Y�HZ@��Ղ����:�3eTp���ﰷQ��;��ۙ��|WYu#}�g
�����wXwV#ˬ|�q	׆ �6VT��_�0��=� Y�p94�/�xo�GF?5������P0�'��6U ��+�lÿ���ڵF�Ġ��j{����9���X ��U6ڮ��P�T��G��(V:]��f9��$=l��{:�G��*i:qq��JE3V`����+��#����M�.��C�n3���f���"�Ih�0��F��t�h��O 7��M�!�w3�W�~��}땂�-��)ּF[�2Dk����OY7��?}h�UQf�M�PI�'��Χ�^zYN�T��}}����6��}|����k��"9U��?lBR��3�c��e�"��P����E)���(J��!�^��H>'(�#Z�IKR���M�#�2b�����,��� �X�7��x��YG-\��4��|)�̈��N&�@���7���n�.Ďo�2�
�?��?e��HX�"#�Xv�.4]Z�!
uǁm
��z>� S��$1�W�%++�(��/�g�������a��y�h�tyk0�^��$6��P���&�zu�t�?��B곸l,s�he�Tb���m����<W�]1�&�@���_�QLy��i���Q�|;;p�̵�75o���j��Ё�f�en�NGFh�l^�6�D�ڜJ9&�5�S=x3�|��N�C��a$I�%��Z��Y&�7��Կ�|8�]�m�$hƍ��Bc��.<��9>�ȭG?�(Y�2�qh�!%�.��C��A��Yu�;v݀�,�����ykdŁ1��a���	��Vkk4�M�!��9߰A6�Q��"(�V�ŏ��$�B���Y�y_TԴ���X��%�Y���ƅ�i��]y�z�D�5Ռ!wg~f�g�Ib���-�� ����"��"�3Zǯz�)�V؝S�D���ծDd�A�t(�v���*j%]a��'��z2�̂p�ҝ����� v4eaky$�o��f���[��w�@�fT���Ce�w(]"լ՚���]r����C\yަ�ews٪�˦	��� �\O�2F���[��%OJ�E��#��缃��Ĉ��a=P�<ћ���De�c��V�-[BM�:����WA�5#����T�g|P�_G�h�����EU,J�Ȯv���A{U��	e20�Ҿ
veD�s������rwO N1��-�ՑTqx^G�p�t-�'��N�+����Rq?'o� .�~F���O�V����u�f\�����崢b�uz^�[}�pL������)�X[�K5]�w��"U��I�|�$�=o�&�G�q��1)�!1�hS�-���\�� �6�}�Dr�ʛі,Q]@KE2�^[�=�\s��Q%��{^X$Ř�� ȩ/_[+<@Dna�~��-nI�P~ ������KD��6�$-�l`�u��� ��j߭����uUV:1��_�&�[�2C�N(��Z���Y����n��d�_���������[U4�Z�'7�~�݂U'�t�eJ�Z����w�v���b��e�ğNݴ��>G�s�����������EɎcE�N�w/霥j���E-ʇ������ ~
�h��<dL���}Z[D4oyW����ȁޠ)�`�
C o{��i2sR&��'�e�/�I=:ɡOP�C�@�AyV���Q#�{�Rk�� gzI'}L���F�ZŶ���BF��ch�1N'��{�H�07云���37R���s��s� �s��`M�X��%;�	��ܽ�4��,f��q*
��:�CI��b���p��9��Kpny��\��Ì9�ۜ%��~�ē��h���2�w!���c��E�O��m$Z"G�5�e0�`#��-X�oC�LGQ8�֘d��.P��ZLZ�&�5��>��y��n��4�U��h�c��)��l���\"��Fk1P����3�܊s���V�7&�q��r�*���b
FV�p���e�
5��g�J�n��$�����]g�����h�Jt�����=Hg���������MͯD�����matQJ�3�(	�G%<M�7����;��zI���΁%�-$���En/��GY��V=�"A���y�Z�>��A��b���Q��a���B�u��ֿ��_���ɢ;T�Mgo=�
�|[�ڢQZ=��Jz rk	R�w�*�qQv�d�`DUb��ɞ��V�M�ˤ�2���(�� �*�|���y��WR(`����^�I�4mM��{��j��k��չ���v�rK��e�Z|���yT�M^Ѱ���V���<yhg=~�O�2�H��)-��DRp����%+o@!�s�ۂO�-$b{A�-n�}�*}^"��V�Q�,��W�Nڠ�?4�쟉�MQ�i3��M(؊E�X�ڮ�<��9j8�&�nd}!F��o*�����j^$ni�v�͈U�e�n��B\�ef�����4���"�>}m��l)#x1ɭJ��[ ���]�'ހEM�+=�RY��:�5�#'�50�����1.F`@H��L�ėRFP�p@��n�B]t�D���v��Ų���I9�$v�9�'��G~��E�S�6������C�Z��~��(1�'%7ն�]�l���{�Q�����p�xxa[V��H�>��-$�������roU$�Pd��W��ꅵ��E�O�+���>��Z�T�o>@�Y�Yme�O�[إ��fr�oT��Z|S���a6�>�wY�,��&�L�o�tc~����L�u��V�=
�L�"n'0'K�]+�5j��Q��*A�vpV��S�w��G���+���K �NT����ݚ�)�W?��Q�HyO��t0�T�B��k�W�\@���dU���v�c�r�pw�n"�U�:��F��P���<X�J����O;5��)�̙�-��y�	^mɻ�0�p.1_@A�1��ά�g��4��S`���8�|���U�O�o�,;`\���q$fb���>�˿3F�&�����6���h�\l�O��v`}t�������^`fW�u�j�2?���8�$ �λ]�0V�s�@������5�b���v�x�W��vk?f4� �;��^�5��[���+a���?o^d�?`�csC3�DtT��PB��@*}��N_��m� �9��_D�X�ȡ��#����aJWX�]Y��w>y��xE�Y�C�G�Cw�@���E��x�����*�`�>FF���À�'q�v��%�D�7�e(�q�-�09�N�j�x��a�#H���Ĳ\^=uX
�g�,�#�K+��Ŋ>[�A���A&,��V��o���2���@���ǲ�Ŵ�GHG����ͦi�w����ʛ=�F:�c�� !���6w/4'Ɇ�ؙ�������\�A����jݳYo� ��7x��$ı�d�0浥�l����Y,�{T���H�0��V����^�"޳4?�U����S��l���>i�q�b)��Ɍ��!�{�*�`21e�*�%Q�	��	O���Y
tb<�vL��g��D�s^�E��q%:��Jqh킽�Oc�6H������Ȣ��e:�w&��3���(�.����D�'U�����/UT�!^�CdOd���Q{��!Z߿1���rĞ.
(u�
չ��E��ǾX�0��ttQ1.K�gL2j�P�����Xsp�-h&~�����X���<��aXT��A@i�uWo���/��v�Mp����=�+�i1��t��X5�#�M��J��� �4T�j��H�S��v�lm��XoXS�YC
W���5���Ƣ��l9,��>qF�����1f/��ݐو�P���it��tg�V����L�S�kVɁ-�����&�s�isz�hNQv?,�vi�.E����@���|ޚ+�ۀ3yU�f>/������2'c��n�����t��[���f�F,���H�K��+���qS���9�@�F� !/'�Y	��n ���]�-qn��ˎd5 <P��c*����/Z!��3��>��+��{�o���0�l�$ǜ{UJ�1���4^��m�~�?��)��	A������	�n���dP�l/�!`�l�|��"�;*�>�4H�E mwI�y��ٔ刈UTq��je�(��V�-�t��\	�r�+�L��7��.h���]��̡�����T#𨙅�j�1<
]-������(�������v�*;�Bl���ݰ��ɒv�})+-`e@cfG�yg��;�
&����r�f:3{�(�;�P�:�P�����f%!_W�L�����$�{��7s)��'Ia�����M4n�����NרS��\1�@`�lƚP͝���6;Р�[;���1�G�tNXMh�U��g�^�W$E4�����C��e����C�>�Y q�]!�4��</�Z%�|zZ,@��fO�S���Y^���}S|��k'˶���Gm��ͳ&�a�����sT;�+|�}�K���7��D�N����K�<�3)�{�e�lЮ8��%'զq�����9���/��8�,J��Wf�^+l"4฿ S��>!���x�ٽ$�0�*��dvo�K�^W^��;��N�ğ�cd�Râ!�<.1Ŧ�+
��B6�Tp�h�N>om��/!2M�Se 'u�j��{��3}�J����fLFЋ����VH7��/�\-�Ϋ2�ӷ@�jN�[���Wi�r5h��p������)��P�����"����������R.�3�C`�_N�Θ�=:a�u&?�/�{]��o��{:��>XԈ3Fb�-��+ �,ǿ��T����	B�Jjj�=������.2����A6v�Wsv���#��Z5G�Ϗ�~J;#h��%���8�\7�t���?�=��`�a؏���d�U���gL�p���1R{�z��g���٢V�u���X���xD,*O|ڱ��lʡ���O��M <��J��y�Y�ݪ�HiO���(Ҧ��7H�js�蕴I&���'y����U��(�� �E����61m.!6�~]W��k&y�d&�^��<�{�W�eАW_��[��Y;���p���Uh��"Y�ƪ{?t�#4�"��S�!�]�M��{��}��j�|c��f�eG��F����IFT~��Nˡ/G�c��go2��%&�2d��(�0�W����ռI'Jų �\4X]'��~"(�����\���Ļ,b�%�lL��g�}�+�*b���8ޠ'���) >��#�;W�Hò$5�6IK���2�SK(Zb�ن�)�آJ�y
�h���R:>�0�� Ƚ�������Z>���ZC��\ŰB�Ɲ�$�4�DU���q�DDr�>"��Wk����ƹ����n��?:�Y�\`|S��k��]�>u�� ���3Hf��8�jA�[Z8��j`
5��W�S6�F0�V_Rӿ�↚%#b^���=��{.�<$�8��iE)�:(�;?z?��?�3%�j�<��� ���yő�r���{~
�����E.�~��;��p�ؤk���g�����G�AT���L\r}4��i!�;MIJje��D����WGV��A�텝�K���m�\����ʴ�}3�D���@���ǹ���0e[���1��L��ݰfp=�`��l�tpp��Q<�W���1���W�}:��/W�`�sD3��d����q~u�o6��w|�t:�|{�.)1�pG& 	&�O��
d�s7�Q?�;�L��c��)g5�P���;f���"���Le,�]�#��R�DV��w��`�V�`����VUku�`B�
�x>Y�<��ѿ���_O���@AN�����}��8B��s��P��(�b�nޅ��h�ݮ����qP�-�fO���1���q�}~7M6�+�e;�zm�U��xr��H .�C���hx���<��9��+�I��;,Wd�	����#��/r.�X^�n����L�|�Ik,�@r�wK���S3x��LC"���~�Oe���9���-0���8ڽ�*�Q�)5;Ym��9�S�?r����+t�od�( Aw7jE�#��U�=R1�=�]շ���	!�{�Q��Ft�,����C$�_R�$�j	U�!��+7�.' �!�1����k����o��A�!�8�l�����B�k�CK��e�l�2�e���N�Vv���Ct�GH�e�@`ԫM[@�;�Gֱ,��#�%򜿲hZ.�Q�f.�F���:¡�w�*T7wN A������[�����t�o���_�dQ�����A�D��zp<�m��o��h���k���dC��m�f'���@��e�&���iU"E���/�y^,b�	�l����3Q�����,��tM
��0{-;��^y��|����p��CHW��a|��zL�z���e���.7�u��r`��%��߹�0��}�4�v3�FT��7�4���s�Sۄ�Г�udG$%�W��5A����#�A�	���"W�q�:h:~n�MDH��2,��a�Ã=�"cd?���RR ��}瘋��_A�o?n��B���32? ��X�x>/N����x�����>�6[���\Oc\��z���<c^�f��꓿����C�U���J<����)y�-'�Aďr�g�Bb1Vw�H����y��{�o�_�!{���#��г�rK!ߞ�����B%��d�C��%��缀]\�x*�À�>T/~Ξ7{hh�c!��ע-d!k�^�P��q��ӯ}�u 5��T�9|�oűu��ZG!킗��<Arҵ�	�XO��\�w��L���FI�3�#�"����Y�����,0'��EƘĺ��<h���e,u4�� #-v�e pB�8�7m@$��Z>�Ƥ�B��c
�
��;�/7�R�l�!��[�A5Rz�);ּc�l����-p���J�0���=��x'����vف�{y�4����n��b#0�.�z$�_�$d��;���k������� ���?h�xI�Xw[��c�#����A�j�>�3":?z�F��T�{?ȷ�i�(#��2��aЎ'��X�˯:��|�M?��8��bfU��~00���yκ�{�|� �3��7�������aU,a���D��uD�°;�l?;�I�&������W���X�vo#o׏=N�ѭ��$�("w����~u�p#�]7S{��.��~���BvqӚYE�Pk������;lٵ/;U'� ��lU���e~:��qK�^��V"�9"�_���Q����H��x��7��x6��<���֥�����l?uC �=�=����ݚ�Mr,f�1�*����v�A�"/�E�z��P����s�y}4O�ψc9F�Y8)�X$t�<�g7>�[|ҿ��[�zY���FɿQu�FK�.MY\�!���ֳd��<L���]���i��2��6������)�-Z��e��3��i_<!�М��0w���u��D �_��%�ǉz�4�Խ"�JT�\>Y��j����:b���p���-��L1�X㔙��m�V�/�I'�� d�A��M�R�	����Ƞe�Z�c3^�O��r��>�h���u��w�y�ެ�N�W���<D�u(�~���:9�t�ñ�S���l:A.r@;̮Hs������O�w�7���s�*kG9�8G�C��_�@�
T`������:g�i���yz_��}Q���I(��"��/e~�;0/�����#�(�a^�H!2-�^�[y�LN�r�xM�\��_2E�<�-3[ ì�ujd�%�o7��T@��vyp�ӡ��`�궭�͜f&�g�Ũ��+�2��]��lު�H.5�v�P_��X�X[}*��+KJ���d5�4�<j(q�g��	L�����|#u�Ȫ������ �|����,2l$��<@�ʛ�2� -A}�߱]�����Y�J(^�du%�{Q�=�]��]}ӽ�ݯξ�QO~�o9�F9pL����	��C>�gH��2R3�}zx�D��S��j;=	Ȓ����/�]I䗨Ǉ,�v�=Q~��4����`�Ԟ }w&}�[i�\t���	��	|�Q�"��[��LM#�ҕ��n��*���$�wIH	�q�6!3gk���JYj�`E�n����"�����ì�������&�\�x���d�����8�h�b���}Ť~�R1�B����d�N�i�Ky��ۊQ=��x�$>O��m�<���p�f
=�s�3X�J5�%?b�ٿ�A�70Lx����)�"	)�8���u]�_�����t��u�9yI�]8:�_&�r���J8GL=���t�1i���K�sI�Y�Em��[��me�U��+
��[vF<�jޕ��!<{�p:#[0�0X�WU54���_�*Ƌ�O���\%
p>�Oj�[��e�����������SLݴ=]T� �}^�[5���c1SCh�#[�y)+2�F'��挹�`D.���������+�+��f�x�  ']��|�+�`1�@e��5]B���U��f��w�&��E};t�ͼ9���a���8���?8P %�9:/�7Tc���It�A1>��~^EC+�0X�,�?�e��#�5qF)�� �r�Ic�~D�"|�&�ݲ�-�ɴ�Ф�3)��F�ys���QlL+�\�=�8`�ܕ���?�����/c�����>fT5���b��	�G"ڃ|b3�m�Y55���M�z�4��Fs�ȜH��(�s�F�6�p�p��z]�&q��|���رhkL0j9h��"�ʠ���Z�H��/q?�-i�|_�`~҂EQZ�WQ�2����v��m~u�=�Xrr~��ܴ���)م&ڹ����6i����Ϗ]�h�n�sx�)�k���xC����{�o�Qէ�6�t��fL���V})vR2�]ǋ�yP>�b��t����o ���|�IE[�@l#��g�����6�8����݃#d�_F2ՠ�����Z@�Z��� ��5���;�S�D-f�&���b���[���i&'�1d�1����vn
��lf���B��2��<1G�[֨�?^�j���-���~L��u3{�/�Q��V�� ����������	wO���U]�C��j��c'{%�?��T���}��R�zR�OQ���\�w-�4������LL��DJ �9i˾���vr��B�4��3��)�ҥ?����|rb�s�*��v�7˃g��n��%�����s2c4�N#�Ig>~�y��i�W�fﱖ{��XKޗ"HK:�LnĻ�Ԗ)�Z/x�`��6�U�WW������tRk�a���vf�����h~�#�*p�<^
���$�:X�q���1�r� ��l0��_���<�rs�at���<�ע�^8�������ªZA���;>ɛ��)���@K���Sm��
6 ;����EH�8��}�jqfi>d��۞�W$?�~�);a�&�[�k>�������V���$�$$>����z�����̩��uY[�4,K�	�+�nhrQ؆���ȭ��T�����(���޵�̗	���&�H�!יg�M�b�O���z�z9��D�7���]�!��R�D�z�`������~��i ��Xo�U'�2� �֣��
���}I"Ͼ
*֨UU�@���/��n�0�	�S��s��V�\�5�YHEL%�m�.��6G���*�
Қ�j�z�}����xҡ�8�p�M�X��4�������d ��}��p�m�D�^F�qv�����ec��"��ɿB��g�"8�q	���x}��r\"�a�Aj��E�G5+�B����VE�i� h���Y�t�X7O��쒼�i�a����j|�áڿ[�#��%%��{��4���.ki�>�5i�y����n�'���21"ݧm_z�!`іg"���]*f�+��]�Ρw��������|�l�
�sX����09�\'����	�E��ܟ^�:�x_S|ZQx&^M�H��t��|��r.|�Z
�V���y	�g�0+SL����+5�����ys�*,�1����$�',�9�p���c	p�;j 'dPP�=s��v���0��L�g�����Ħ	Ì�]�|�u|N�k�O Բs���΃� V�7Q�b]�������!2�	Q"�)�ӝ(�c�)o{�@��:*���r���[OHv�����U��E�P���,��v�6�>�Y,�eϱ4٭���,J�����ao !���Я�����$G?,�F������d�b~�L�H�4��,";;��M���a�}�?�@��Q��p�t���������7���mg4�����QQ�FRT4��a]�x>�-%����ՓN�=���F�bWU��r�����Y�rU9e�-��+����`>�F��C|�_M��"�N��;<���l ��_�E���n�#��R�5&��^�'���k���� &���zi�
^���Z{�7�s�9��/,�(L�������w�Q����}�[��=�6;�AÞ����g#Ƌ���3^�?���ޏ�|�¶b�hN�k`�o����1�y�/���ET������J�.]6��h�Яʀ��
`,7b߁���>q�n�?��U���ߤ@�����}@�\�g2��K��#!�k�7�%eLj8��rejx�%�[�NV��k�?7�S�&\��U�C�3C"�@Oj���wg����{h��Y
Oj��+j�O��t�Z������2�5Do�c�6�?$���ӏ�ݴh���R�gu�6~���K��E�O�W�Z���[â��K���	x q=�
8@/|s�&Y㏿���~�Vv[Bw95���7�KE�n�kT1�*ࣷ������x������^VCؖ;�X�w21�T���f�ˬRB5]�9-�c����1݅/�z �q%1[+�k��	5�2E�C�A�imSq���X��pj���I�+�P��gu�����g�bL����cQ��fｨ�uF��ޥ䀈w��qyz�(:��x,�N�7F�L�U�����ZIتjn��m��j��"��>-�
��trSQ[C�ק�q���v�8!���?l���RY��3f#�
L��ͦڸl����ڰ���V�pv�^��"ecMQwZx��f�#�Â[F���Bx����/�2�ְX�2���l��Dҝ�5	�	��f��Pn�OJ�:Bw�Z�?�̙(�D#�h�$�Q�Ms
��d[IK��L秂5�a�;�^��W��������`0·8mG�5����Zj�?u�\qT(�͗z��V���?�<�`���+�IX�DS�`��h��*r�u�γ9��XP�sY,��8O9NX���L��,	_ؐ&�)R#;&5�%��dDـ�9%1��M����.��q~E#Vze��7;�5�;��_��IY�����&7P�8\��i���'����W�_�#"t�K�
b�вl"�ڄ�J���}��K�]'&9����h]���m����}'Dh�3�
�aO���-)N�C�rA��@�CS�5M'���\*��-r��v�N�K��9) ��C}�KW�7�֮�� �a�i�A������:�Z��Vs{{Y_��SB��O?ƽiý�������2�&�'{�ɜ�n���9	=쩙�b���\9�_�í��dqUlG�q��PZ��9l©[����JV]�-�ҏ�.� �+���A�=	P{ �k�e{g#z�c@1?�����Ƹ1w ��khyJ��c��Q���N���|�p|H	������:Z���vBK������e�$pX�������pI�,�\۫�į���';B�bjAį�[�S����!v���`�
ѳ r<�'���%ek�{�0�e��%ŵLУ���7��̒D�	�_ ��p�˃�%G��64�Ց���I�}��`	��	����	�g�#� G���u��8��=C%'�N��r�si2�ux+0�0/Î���H���&�-�X-���C<v����)���O,@���ux���G���ڢ-D2Ϸ�����c���
F]O����k�1�ʇ^<%k>z�1�oߜPZx��Pץf�?B����8[~�5P�w����\�F��c�8߶*z��i -=$CF���W���&�W�8P����!��w�3ڐ���|ޮ�5lp�`���߄MR=��w�
<A���>e�D��o��.�r4�����ƃ�݂�`����x(�_�I�S�1DTVR蜁H#�!j��ʒI�k+�+O�!�0�d�: �3�z:��%��C�T����2��Q����HF�|k��Z���Tc؉V�Q1���I�m��m��Ij���fTCG�|��!����A�x��J�Fƃ����ˬ�%�{4�({�Xmk�u����1$��	70��f��KO��ڝ��6�m�}��HR��;��Th7$Gbj�̱/o��dr?iVܒT�5T�?����y�5��e������\����ي)h`�՛��Fl�hɛ�[�˜0{����{�_��[�������0�4�-�"�`�܇gf��M^�4���Zdd��-�"�u��
������#,F�f0�s��O��hssia�n��m8ɐ��[����A;-ࢿ�0lʼ���em�j<ʻd��f����i�t}f?]g�E}����za�n<�s�nD-�	Ѥ��Ӡ�f��z�z�O��Mפ̠�Ӹe�|s��������	�_�X.G'�M2�F�����zK�a�z���c��A��rAe�x���� ���ph���!�+8�Ҏd��ˠ�~��P�~�0Y�+��Ǔr,I�ŭ��J�pm��&E)�\��2���rd�f���B�3�+mW�M��~�Tq-N�e��;�i�Q 0�=:	I�6�}����TJC@��}\2�	+��>����XHs�J�y4�k׵z�=�G"��=F9�<J�z�۱����Y�`!q�ɧ$�)B�j��)+¿��[L�?pD��� <��E�}P�$<�y�>����1�ZS�hbJ�?.�*q_�+����7����8�����t�T����a�:')�Z��K�ƀ�* î D�P�j��>�،�ks�� ��~�F�*�z����شi��Z+4������% xș�-�	¯�()��J
ǧ���T��ubL埌�gKf�c�6��, T��1�»'�zX��q���i�D�8�e��Z��C�6��7�� ?o���������$D��"�u1���"�^����/����?Lǣ]� ��5{����;��؎�
��ۉ,�t�nF�X�yͲ��J��tK2����7���X�wg�He��p³�֯��
��k�!k޾В���SZ7'��4�-:T9�H䋺�3�Po�4*��iy�b���I1P�Y��#O��o
:N���ه�M+��q������؟s���[�����3Y�jM� å�]$�bw1��fh/d��R�� ˕tQ#�f�kՒ-]�v|�~�:�E9_��#3�
;�?���x���rDC�>01����Gl�`�{����f3U?ʮ��x��ei���߆8�lS������g1+�B�3�_��L�E;�\��ru+��bL�o�[�c7��g�l�'��Jaʆ׸�����A%��Ҳ|�ig���woXaj&�1��$�a� D��_����㲣�zYѝ$# #(o:ް�#��s�ě����{	��'��z�t��`˽�r�tm������2j��TJu��7�'�\�	ʾ+!���A�׮.����`*�_�`(c�Ȓ�a���Tj�ٕ���'iNz!��� ���*4�vRC�,d\/_/��HG��n.=���J3�}s�cBLx���/�(������q��/ݜkB48����ܩ�6�V�����~8�_�"�tB���_��줎�I]8�d��;��Y��;���A���`�����6y��iY$�d�/���9}��>��l�Ɗ���k3F"������Ư���dl��w��z�w���@�%�!�͐J���>t �/CS���=�l����\���U�L������I�Z�|�Y�WF�� gf��Q����U���(b��ͱ9��޺��h�<}i|���c�AF<�� !����� ���u����D��\���A�Uy�,��'��@]`�q��-[�Z w�^|C�E�P|cc�H^���!l��*ϩ9F�v���:���̊1���b�{���	�k6P>�,�����؄����#�*�i!�Gr�v"zf�t��b�X���qA�F�{�)B󰮋é :��U�a$D<�@�ew�[1�WȒ]� ������C���R2�nޗ7,v�L��"L��cZ"�v��Z����>^�#^�Pu<1}����{=�H�������%�-��!%���}�r�����Fy��.� �]*���&��v*���}��BI%~0�P�h�h�ܺ8���r�Z����)�
�� �"F�ռ���e�tךg	ي�Uh�GsP���`������uF��%�O6�n�ª��<e�����,fzw[����r��4T)ˋN6`\#� (Ji������܍�i{!������b�����K�7�W���I����H�����#���g�UU1�lt��ti��H���g4�:ƫM��P۞��H�o*X�!bn#kk<�*�e>����^��.$cr��ı�Z2<@9���^	sL����͞��+	���_�#�V�|��Ǣ���
�){	~����;��h��MJ�O�W�{bK�,�MB�]*k�%ژ3g9.!�oW�&�t�����iC�v��HI��Pw#>Ԡƻ���!7�e��`�d�f�#��c,��[b�%�ѝI9�N�fH̥~R%K(��mÛ/.��S���L�/9_�-j��3�A�ij~����k%��*�J�Yhi����bTS�?ܫ�e%,~O�A���~!�ך)%ߠ�lĢ�ls_=E>~D�q���Մp5͢�Nq5B�`_h�}�iMi]�<���Պ^O�dū��)�B��ϩ \�DE����հ5��n>����������;�3���ZY��?h{a
��;�y�!6�)szD�W=�\Ʌ����=&"_C\7��B/,�U`�	=e�zu����ּ?�Wt]�J�f�"g����u��ހ(rvNxrM48YR�v��2u�=�	Q��oP}��L��&�r����蜳~��W�|�h$�|`k�5�%g��t��n���h�R�t�+mOH��L��E��³�:qS����^}e�M�!aj��ۨ{���2v(�j<���ȅ��İ9攋�c��:!҄������������r��!�\W�I3���#�h�v���z��*}\��y�i�X�8�*�y���7�a�M�;���GpX�T�s�G�^'�2 Dp���|a����B'�MK�(�!���sr��A������o{M^'��Յ%t]�"iѶ��ò�����=�����O��#Z�6�R������O�z�Xl�W�8�b�u�6���S���?Q�.�b�xq��ѥ!���-k���U`��v�a�������5��$��^�u_|�}(��ʺ)��i�UX�2&�zM_���s�B�.7���@�FH���35��7Ԑ�	B��HP�bo��?\����,��n!!�Z����ͦ
������,�Y�F����K����H�~n�#������qZ�ڨ'Cڷ�D�&˰5p㒘�ɸ����Bס:u5��l`�.p��\8��KGN
DqKm��Ԭ.��:�%��8��g��»�V���I�{\|{��K�S�̯6#��JM���]��?���Nέ���鬏)MJ�O_�a����kÁ����"TύK�YPy�����4g�Ǔ����\_|���u{�F���#��~7� ?O�`�l�_�z<[�\����mѺћSY���oZ��q��c~d)*{��t�;a֬�yAj2���F6,Ñ�4%L"�??��H!�>�,]\�,,�?8�Ǘ���|�<u�`�o���xO|]�����J��@���i�4�u��
?b
�[دZ�Csf�
Y��p�tK�����<�v�����d���<,R�i��3]
�˪X�2&"�Z��#x�B��oS~�R$~B�v�.^�%<�sAm���Xl�K*{���.�������]jV9,�sQCE�q�����R����J~^���[�>���]-S=@.I���5��e�"�#����p��C�^�R�$L�@�wT�K6
�	šg��D�`��T�sb�˔/h�(� �����?Ī#�<�=$uK��W	��L�����]�=##��r㋶�8l�HЭ���Dv��=S��(O�7�����L��tXR�X���P���- u�ŉ�3����&&D���L�,�l!p$���ɥ�z�T���A����+*R]��x�0��&�/���: ��C��B�����Q�*f��7�R���5\��=�8P-~]�q�I}�L�$���.������@|