��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%��F���/��f{��$����	��`<^t��r��%��	���;�5C���(�� K�@ӟd�jT�1�������j�l!2�T�mf�v�}G�^M.F�j�D�U>��j��I��vT�]�M'�����z�E��=!s�=b�7�/gB���X�U���D�� J�~�]���e�R-F�o�t��1(�ɟ��	D�]x*Q�*�W��߻g,D{k��qhi����YJ�nC߱�l�ſ8�D�l��@��(!��Ll0���R�"�{l�����9�a&0���1ij~`�3���3��8�NP�xTꠑ����~��я4�Ҷ}��7nV�Qo�Ƴ�J�&�5�������:�rW1e��g@�ju�d����A �S��Nm;��GN�������rO\٣7F��9s͆� ��t�B�l�q3��P_��z�[�{�t'�xu�s�4������]H'��V(<Yܝ����h�Z�R5��h���;�DeM�*mg �$6|�	�è,�ӹ���ђ��nDX0�@폂j1;h��:�e|ڟ�p���V�#T5��6���x͂�<E�hxF��N�rߏt��@(�Ard��Z�s�@����i����q)���r�z�N4�f���b�3���p=�=�Ś��/�<e�w�����RB{gq��կ�EF���88�	6�a��;:�m�m| ��N�~�~=.���0�kq��-j^9���,L !ӄ���a:��8xLk+��x1�fN�p��^��q!@�*���d��u3��(��bm�9���Q��T� �1�'vp$��?��f'��zܺ�J�|��e��"�ay�ܪ9)�������@͘/ؾb̧�����!����o�-uGz�=�X�DOq00V�\�H��݌�p��4]0�o��0{��`���}���,PIHR��|߿	�֑�)���[����N;M:N�J�LKm#����@\��>�V�T!��q1�V�
�����6�у)�`��ڈԥ�e���"��q�(�ii�t'P�ׁ�5�Z��I���iW�²�7��tFh׍Eeu��h��p*�v�&�4YX_1�e��3Ŗ���P�ō�P��ᜱaX$�Mh�]�!�t�vs��&%���Q� ��}��d��ncN�R�FB��HN���+��j|I�̺��&�B/Ѿ�Dj5�r����6.�=s�aԜ��a��H_�]�S��`��U���جX���'�ϕ�K>/�_RP�)܎�(�@{���^W_2n�(��=�Mg�p$ޱ���~�Wz�}97>1�ٞ����I�	�K� ����$^f�zI��Y��׷)��z�:�G�R:7���<��;�#������;�|wz�0.�clN�A7�h�p�2U�'����ju򩪤S\<j��yսWG��9��>��5�,F�$ήgś��\K�[������QYNt%蝬h���r�6/Y8&�eĉ�N�1`:�i<�Sj\Ǽ�5M�a[�L)��
��	p2+��P�t\+������N�_�?���rCeJ���r��M��^Z���螷`��=��G�aܼI���Ռle҈rJ/�B��BD����"S��cV��q#��~��\(#8����+��-͊�n*���b��px�v�3,}��xD0�ԝ�Z=	8L�,����}�1jу�<-ʦ͒�s���ϸ#ޒc�~��%�ڧ7��T�'���9�v���&�:�x��qm,',�ܟMu�ٝd��'y"�xI1f��d��&Qo
V��&j�ƴ��P��́�,jK�1�s����pWŃʹ���a��{�K�v�e�E��8v�o�C���v̝?C�V���0xKQ��T1�����B���I�ͼ�	ڤK�������ϋŖ`X����$����F��q�}�Q?�65#|nG�qާ�q�cGN�%c��ܒ]C	�	;/��n����#�x��Yuܭ�����оž]!c��λ��=�3)6��Đ-ŗB ϣ�2P��K#�y�"��FL΄�W�?���G�_ƪ��}l(����^7u��=����	_`��R��r�<$)j�| �D���|����}p��)���n��7C��]b����Wf 8Ӿ��|�l�ΐ�޾�FA	��
����/�Ⱥ�C�.�����&�D�{�Gٷ��m�"O J���E�%�n��-)CZ4N��+}#+@�o��s�05��ء��(F-��)2;Ka艹	v�P��
ї>����mZ���9��L��dȋ�=�5�e�ʝ�|�s(�#N�ɣ��uA���P{)T�З���9 �������'#\�~�n6
5B갍3.�Fє���{���#4o�>\C,?+]�&'����jSQ��`���F��z:#͆2D�S�d�.�kӝ�C6�և'3ftt�Uju'y@&�)������^��w++I�o�M;NJ^�?U�f^��QsS[�#�B��Q��)�T��M)�]��܌s?n�ݻBY=1�H |sK��IE�?�R�����N.�(*<�h�뀏^�RWG;�\�U���jA����?�~EZ$��1OǄ������ZЯ]��ԋjB�Y�O���Ú_<\\���Ow�7�Lם�����X�I�Eʤ��� H����ޯ�ٗ��39DK�"*��鋨�ױ6_)�o&�v
����@�)]E&S��1h;�e ���@!R�W������yU3=b^"M���m����زw�CfKG��U)wD��̔�����Ӄ�5H�t�/7Ȯ��n�yĴ� �����f��@��;6�����9�4���&~7�����Ut���F{�uK����1�'H��F��
�7ƏH��8�D�W��3s�8cC׿���蔉�k��.�S&�<�̢����==2����{�#�<ߒP���
��v��TƮ�n��t����B!�N��,�je��t��@��{��q�ӊY����^�&;ĆX�z���qP�Q��:Q?����>�ey�X&I�c(��/�#2
\�I�k?�т���j��n�-ՈKH ���d������
��J�� ��e �7
�����o��{[�.+�2� 30"�� ���_�R�k�W7\�Lf�n�����}�%9�m~�O���
r4±�NHJ��:!(�����
�I�Ed`�x�+��U�)�DU��Ώ8� �/�T�,��Om	@�?��d��C������Ł�ؕ���*��6�+��:>�@�3z!���J����.� v;����t�����W��c�ѩHz"A�B��z�� �H��"Ej+e��@�G����U�l;����*s�2x�	K�7rrjF�qi"���C�Ν��"�w��ah�hh��|�+�����Yl�%z��wV�-�K�:mr�����-���E'Spj�dp�� ���i�}�x5�P����`���	��g�]N�3xc�-���S�-�.��P4zr���5�X+�i$axvU�W��L��bZ��S��H��(�'��ɼ��L_� y/�t�-��)z���.���9������9D�H�J��/�B	��1��	\��J���HM翠��Q�G�}����z��C]?/����e�Igj�bC�Fh���]0,^b�)3����6�/X��y�Ψw��c�<�(�f��QT�p���+%� 7�y! �{����� K�ѝhg�w�W����7��42�.'}�=�~x��IGR��^�cQtP-)ǵÄ�gkmzS��,���S���LX`*�j�A�/�Y���J�{]�a���H
~�d QhY5�QA=qX�k����_ۼº�P�VVS�� �%��S�r<��,����~)wjU	(�f�5��v�iQ���>����H �e�ҕc�@R0%�Ps������`z��b�Lt��V])U�]�����|����B�%ƞِ}2/�ښ&�E-/M�O�1V�U836g��0��۞Hu�y8�^uH}.o�i���㐻����з�yC�vk�ڔP��0!ce��:�8#��||C�]|��q�������{9��E�r�$C�ʆ�\n�k�:�m�i�ŔL��~����6ք���%��<ٰ"����|~��m������v(���@<~8�1ĳ�$��))��S9��[y��Ph���Z���,!��B?�K����T2�|�C�`����S�P`��t#����kD�bT���A�m,R�3��A��nr�(�ч�eN�c���ㅌG�{z�cMaM�����tO���e�R��5�_�m����K�1�����ݲ�J�(�R[y�X�����xG��V��Z_�%3��F3m�����Q���+*n����:z s8s[x���Ȼ3g�l��#K�y�A�� ̖��Aw��[g\p�,�+[��dƆ�����y~AC��t�pD.��\i���]R��>1Kg��`��Q�o�w�s���<aգQ���ؙ>d'��w�XL���h����d�ƶ�3jq�\����,qJ�/ն��y{���Uy�bN.��5�����=>I�I�[�g0b����Ā�@��3��������f}}�R)����,X!�����41����|ō\F���p+*Z8l�Ls�&H��@t���6�W�-Ç�ޮ�~?��D�L�P��^�t�7��o
����pf�Mô�1�I-�X���N�QxY��~�0wz>7&������V��X�@;�{*f8�y���l����a��(�������k"<Z�U��D�rA���$x����Y&����_B�$O�(=�	�W~�>�5�DV�`R���9^���6B[c|hҧJE��`P��\u�+�.L
���h1���*�D�>��^K- `^(���fE�!	�)�Ł���ԕp��IgP�
����R��B#�kr]���S�������������:��l�����1�zF��'%�˕�E�
���jϛժ�W	�9��KŻ�8C	���h�21&�x9�7�M�g��b���_M�����w2����:��o泷��L�>�Q�ڻ��@o�$�HU��N�����66Ӑ�V򘿜7��|���h�J�jc�/����=fOW�D�7�SI]�D.z$�� \�))9jځ���U�')�P���]ό!#`�'ۭ�CdK]�y�	j����s���x+�N6o�&��s��� ������ʌ1-�c�������9A�:�T��c������L��m�	j�B /N�A��1�a�$�?*��Q�{d	��X���ֳ��V-������WJ��pZ|��6jo� <���x�D@�~�=(���Y���lE�u��lf[0�L�:
���33(�%�_�$��\^���W�Ҧ���N�����all��v��pmdAӈ�er �f'zΈ	MP��]���躮��X�n#U�I����Nf�BN�A_�^������zܡ���h�\Aj�4^%�C
�n�]��mv�@�y�O����*�ݏ0�,܇�����&w�Z��'	�nxD\�5��|�p1X��Q��W�~Z�:d����	�d��><H��V��s�b-fJV_���!g`���.�^���� ��|Ҿ+�"�£ڞ�����v���SX`�.�g�μ��7p�h
�M�<�k��������z���7���)9�<b-0h	��c,/��@���� "t䅦@��Ww(D9��5ᰬ/��e'��$b������=.�v�#�W� fk��ڛ/@kS8Ǳ͕r�����q
[�����Ï������ɲ^����{T�&���A��`�0�giCl\����+���\��<8*�@1��Zն�<�y����MhȫY�ek�e�o%���	����D�>�n�0	�N\�A>��n8�P"w+3��z���0_��\��r�3�כ�3��_���0Į�x�R/9�~�Q�(�y=�"��(��2S��zq��ɢ��_17D���H��m�C~#ٸxk�%�js<_~���OXP��f�>h�����[���I��
�}�DA��&옟0�*���aB&�d�eN�����G��>�)_"<���$@{�?���ul��B��9���;؝���U�j�*p�'����z;��	ŤJ�X���9�7J\�\�	�i�k�>o��ʊED,4/V���Fg���
����7��/;|A5ܦr��h��W1�>�c�ɾc&a�2�:�}ۑ�y�8�L�0����n����i<E�OI�8��G��g���ۄY�	^�t��kVI9.�H(�"�ȡt����_�T
�� ���6F�VK*�E7��=��~�x
S�=�j��e`gC��-M#���M���k���?V2����kh�Sb!�~`X��t�|�MC�>�B�E�s��޺mZ�|��%��8�>C]՜ �����$j��������|�l`�:o&�����
�����k>����a ��8`-/Y�˵��r̖b�%�w