��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F������gm^��,�����ao3�_8}���(�{��55���z�[.C=*�.%��]�2T����!�|e���s4�7���a�K ���z���;��l��|&���-�5v�'�#th�$Ψ��P�7|���ɹ�o--�ע	��M+ξr�-��H_:W)Ԡ6w�d,�;����<�5?FT��֛K�m�@�y`"�V�N�����2c�@Əhn�ߡ,���.w�#��[�WZ+Z�;D1�P�����#9�(n.�	�_%��֚��	�;�)��l�>\nkY���@�#MZ��g�� �(��x��,�j���E%D��K:5��,⇓�s"e&a�tZ(f����oEJ\�,px덖Yˮ�/ ��;����_]�ws\��RV5c��/���Qw�+o��C2#P�/�:��?����_y�֒�+��3bv�7E��$Z�2)�H���u�|�BoXoãb�(�/x�A�O !�KV�SB��"�̨H+��현�4�i�tO���x�U^�R��GD>]�5)�9)���;���q"��(�ϫ��/�$��0��DF��j$S �c��^�W �Ӳ*0�m�Q�:n7�8����z���&��m�L��	 ��X(I�B�@R 3H8�Đ4������eOC��D��+yW�yF�nQ�u��a�5�9uv?W\�/r-a�4��U�W.��|��*(W�d�SBz
��Ԥp�<��̼z�{��v]|�%J-�����c����j$k��+ty��FI0��ʪv6-��D��eO2���p�/x���G֩��50]d$�J1�5�l׾�ڒ�=^Ƨ��I�EC�Ƌ�0W��ю����)��c�w@X�B0�r4��T��Ym���&P�T£�{��-sZҺ�Ds�.A��2��[� b�##w��ԕ3"v_g����ӔGl�6\M!�1���Ԭ���7�`�BJ������옩H�ۯn�yo^�&�S���FZ]p2��g�ջ�,����]씉G�;5+�,Z��W�Eˇ�Tl�ov9�"R��@M
���H��}f'�F�"|]��bJ�o]����0��!޾�}�D1�Q#�1Մ�^a��&m�Y"�|1jv�4|e2s���eg #��z���F��դ'
yOվM�]y�c�sô˅�ތ�b*�*��S�F�b�8j?$�������+�4��utg�S*�i �Z�z-�pl�6kL�l>�ZB�n1�.�x+��IE��=<��a:����CO'��c��̢����R�<3}V����$��>�Ll+v%���+������}Y ����2  �l�6+�8
���Y�	��A�B����mc��:�#>�S� �y�X�޿j���H�"��.���ؼɴ��l��$�}�펖	FY�ܘ�-���"�߯�xNEvi��K��~k��sN�R%�j2 BtC0�7͍��Z��}<W�XY�\��`Ķ �d�8�DB��OJ�oЯ)bV�w'����l�&'��b���&�(e�'�;�n��3,1��w�x�`BL�VWjRӑݨ�ƪ�.�6"OsyP xu��/�(:�^��%h_�ʆ��0�U�@�TO\���0��G�D����0��)�D��6ó�^g�'SN����4������(T[>Zx�#@n?��)��4�'h�S(H���'��ڱ��5�V<*qp�n1O �t�ݢU�x��zyj��LB��-7��Z�I�!�8����)�R�Ah:��Zp%�5ѫ�bs�:�g�{Rʧ��!����M��F��C�����gS{f0�Y��(��B�vwD��?&���'iН��
�T��,�+�K�cN�趐�N[��|@J�5>�"��T�/�vן5+9�����lۄ��a�A��Z�Q�GԃXJ�S��ϱ�(��$�/� !̔dwV,�Rdpx�Q@���X���%���Ѩ�;�$Y�!:��5kW+{Y���X�G�z��6z���ba�c�-\��oZ��a��Z&��;.@�3)��ˀ����~�����:��W��b��"��������vG��lx� a�CA�-F�I��r��O/	�φF�:g:^��w7`���(�U�����.ú���Sάw��{�+	���2���>ŦK�+�D(�%��RRb1c��(l0����!
?0}��>x2Q�ʸ�6�2�����.��T�M���S�� �������%����:P�f%��mnn��Dm�n%N�w
�cM����_�WJ������Y�G%Ih��|�|��P�>]�OA��An�&S�����Hf�zs�ɉD��VC�ښ0f9�VT^�{p˂�xj�z�ر��+/G�B�����Z`�������2�Хݯ)�K&�N�q����z����p�T�r��8K�K����wy�^��eko��&GBr���M "	�u�@��K�s
�)i�d�>t2�7�$�mNH�ޟ�O%b��YkvuP�H�<�P�*f��&�r%�H)y��e<�e_�Kl���Ie{��J�:��Ӕ5��")�̏6%�F}�.�0�ep<]��B��U=��(��c��Ax�`��F���㍙�e�y�'��@N��� Z���ˌ�: P@�WȮ�XK��{Y���7D����2D��*�|��$��)0��X��+t౜�{��Um�p�=�;�h�{-��!���£����|s���\ꚠ��������b�
�6���+A�czu��I�c���{C͏�,{Ʀ�������'���]33eH�=�n��:^qTh���4k��	`��Q����WSs���Qf���u9�0P��f]J�G��(#�I0�(��s(U�0��^��
�(��ɷ�Y��Vh2.����2��I�S�F���>��N<Pg2k ��)X9�׋;Y���(.�,"���05���h��������9釹zp����N�����Yw_F�g��*;ĨR�Tj�६�Hx�C�8�������	e��3�Ώ�h,��Vk+p>Cb����������ꏒYX$�혘�k挆�5鵤u�@�#��� 3a&�S��1��Db�>l�M4�>�&�$��c�/L�R)0d�t��Ј�WZ�Ҙ���F=Պ�r�LƳ>x��*&&S�ܓe'����#��Y��D���.TnS<��|��n8R/tw-����i�:b���W)��������9���F��Y�Hr�B%�(��
M���k��[�2K�����`[1g�щ��F|В�i���=ʵ)B�x�����^�Z�C�<bnM�b�>0KȤ�;�c��"�h��T�-2���">�7?��+a�
��I�I{�'�lR*�Ψ���%����-����e���"��$���|��%��)������M5�{C���Ñ�K��5�����\6� ���ڛ��&@��Ai��/�Y&��m��Č )�������'�of�؜����i8.*��T��jF���ς�`n�9����l.��B�α�:ǧ
b{����!-��Xțf�/>�)L�8/����o�R؞�}��=U�{���%E�j��v�m��Ŏ�@*���Q�J婤� �*ID�R�
!�����*��Ƙ�C�����@"H������~` �+�^��^�<G�9峙SôZ�"�SRA��>t/89�mZ#����Ǭ1M: Se���5K_�~������qi-[���^��p}8��)a�����߮��U�C�'���
�b�ݮ�e�_W�����bw;�4������9�g>Lt����I�!uￒ��S����AЛ�'\ky=�HO�Hf|�8>2���YR�0ADm��+����j[w�r��UtG" I�uU���94*�%g(|Z�àO�TM�vch�H�]� U���ֶ=��O���$�^��$��F̶�����Q�]���R"�㫓�=�6l�����<u]��w��w��r*���BYR�ȌT��،�˪�l*� �<�����E����\^"�(�Ê�X�4Ŝ��>�\��XJVUP{� �՗xP	�Ӑ7��3J��Ee�)��MGs���e�����;^��@lA	X�>=_�v/G�YX�r����ҡo@;�󢹡/���|�>���[�^H�)���3k�.���-\�'��r9Iu�nJcm�'R<tqw�#ܬy�Zӯ�L8�G.TA��yx@�c:a�G�c�G�p�=oȕQ��Iqy=�R���T*����U;�ƣ�^�u؅������y��������K��ka�b#�W�3���E����.��YM,F�j[o���8qΘ\AG�R��^�l��t�3M���/:40��	�Qpd��{��h.7ё�@}�+ h��z�����tZoJx7q��0��Ui������ܝ\Ɍ*Z�	��˘�ߞ��!}�V���a0<!o����� �v�0)��
���h���g�ZhN2bn���2>@W�y�� ��]��|�ic�.(��dD��#_�U���(Rˬ>�rd���7���qR�b6�y�j��C�iaן~:��7;m��p6ʖ�8}v?���ݻ��"wX�3W��� p�_��?��?S�k���geE�����_6���wF�zK�0��V�򤠬
����=V(������ӈ�\��9e�,R�	���cO����N�����tѰ�$j�#7��<1pC�B�[0�+���+5���X���C��{�o��	�I�)���R<#{�{8�rCO�򅳁گ�F����f���WR�"�C�}��г��lfX� }��Q��Ҹe��� �jK�`�֯t�(���4����{�\U���bz=�Z����<��Τ-	y��2{�����C�����Kq�{�M�t� �j����jy��i��G`�����F��n�z����跚�ͨc�����_�ݵ"�o�
�;��_S�xq�m��AV��yN�	NƇ�-%ր�iw�9-�P}X���Y��̑Q�0���gâ@�HEY��l:%�I�`�K/�o/�=E/�Y|>�d4m0�x���x^�'R"Ĉ9�K�VlY���oN�>y�e����}P���c�QnF9�4��͖A%C�����{� T�?�o��s`����]�at��:R�7�;�;a+ghL��~���	�B e�5�h�#����ŷ3DCj�KX�^�o�ԉLMA��ik��-�u��V4�guI�;�cNx dP`DNI����T���G�yu��@)d������qXn����mDrU�jgZ�h���LG�3}�G��_T�x�u������=�jAM=���x��%��U-o��n�;��s�E��}��"Y0W����R���z�)���SGu\:\��Qen��`��B,�#a)~i(d�1N|�3��3��a`�c���������3:�Ei��^^U�B�c3i�H��2������e�c�OPH,��+�Y	�cOc��c��٩�����'��0�k�Q_E}Ćϟϓ������Co��"�@؟$=C��C*��)�G6��R�9�G+��$�?�=���Ėdq��x���%�m+
�� ��1���y��z�O%p�Z�2�>�%%��7����ٕSW�4l̯^@k@H_9�)�H	M��M��s�t�J��ڒ�-ݻ}���������o�ȻP^�����{EnzZ�6a�����)��D_$�=�o���1����y��D��������z�j�IםDIj"��p
���ݧ1�H�0���ϣ�hFn�u�I>:��i�i���� 5����YE5�X�閙�;�$�T1p�-R����'����%���U�>/��N��>õ��(�n� б?�Z� ���	�ĳ�3h&���-UN(@��Z��M��9�͏z��> �kT����:;�Jt�ഠ�q.��w�Qt���+�.�6�\�gBk%�����w�pR���Yt��ԇx��]^�Ż:�j�a��������}b*�$5[M)q��C�MG�g��)�?K�C6�i�op6��K/����2+ѪH<�G[yj����1?�4�zS\�w'_'y�E���h,��vd��r9����~eYw�l���s�9f����?
��^��|ոO�A��a9�3��ū�i�h�m����VⰍ�s��%�I�*���<�I�� T�v��U�x�*�J�3%�J�nՔoV��oӾ�A�)]Q*�m��'7�7<�2n�K�o� �[����ԕ@n�n� c�
s���V =���2%�+@B�w����~W�7.��+(sn=�o��S�-�b�a�b0���?�-yO�e�����Εfp�.���E)�_�r폃���b⢏bݙ��E��Lő�E�׻ˇCu7�t�)I���X���
cV�F�%�̔�WF���E'�ᦅ!
��b4�mߋX[���M����W��B��=�����<'-�n��h�C����Ra��u[^�4V,WfǌH�3|w�!���&�1.��v|��GLUZ��̔Y����O.�����6Ǟ]|�i+��' �]ӥEVh��M}�������"]~�R�E.�zoP�����a
l�+,𹝺���~�'�NyM9M)�Rх���ǃX�=\���~͸k
j2����embo�x , k��#2n�J����v��}����+$Uk�^�*��x�#�=�C`�*"�u�'�9s qM�y���=�H��1�n�Sk^[�N�����zc^_F���Od���U$^�o�u���X���W:��N��ԁ��[ZG�f� �7U�/�PDL��5�D�%,�ύ5�7~"�9{-�D��Ҁdj��%㯤$��E�~���;��Mvm���t \�h��G����=�(05�z%5�P�����>3�v���@�H
We{v���BA�sr����<ʑ�B����ŭ8�Q}%���Z2�kT$����GP����Y��[���?]�a=�8����槀��0�F�69>=68`���M��F�B��h5��k�a,G�L?I�گ*�+dd��d&�L�T��ۯV���kH�]΃�O����Ԉ�D����B��࢓s#�d�9��9)eR*�%;aM� ���!��-i�P��tb>���������.:�m��s<&L�B��-��6�$^:i�)��hq��sɖ�"�%���oW���xՇ��������R��4ῆ�7�W@�r����=M&1��>}e��>��?";k�|���N�E���!)%
W?�2;�$��K��/<�����(Ψь>�8nچwn�pvI�fom�QH���}�z�5"���gX	|q���F�x�goI��OӯL訅 1��� ��t}�vR1�	�'��������F���u�&�����
8�����W�aì0Ri\��4 d�+����cs�4X�X��0mx,�X��俩��q��m�j$����W0i���a���HB���N�����J�d�����}d�o�XIJ��{]��ƚ��E ��q�d��ku��Q��r��A膯�d�����^�3P�]0��ۍ�д�?����L?�s���u�� j�m�\gS�&T	6�ϳĞ�lbd�:��v�-����]��ND��n$Y77����-N��ԅ�CWhe�0��dG�蜆�Q��G�!w�oz�?�鱔�@1�I��)���rkm��EH��;,-+2Su'9O��r���Fi}:)���ğ�9��^[+�2y��v ���.�����4�#
5��GE\�*�b@A��б�����'NxB�5��|����=��!`���H ��l��%��9EEY�C�=R�%�߇/�~���ɿ��@.f�V�z�ԫNM#N��.y�﷮m�J���*�M����ѭ�0��P�ݕ�S�gBh���)#��a��
0�P^Yx��R��P3hj>��`78��@*C�#����Z��cL)����[R��7Z�)(��I���i��P��f�e�^z�m/�CU��	ܾ�qs�B6�m(+����>��>�\+�v�4{���RI���:�z�ݼ�r-���աQ����g��6t긗9N@��e���w����3I��-<{����b���3�7�����a�#3��\�oH�0Ig&���wNJ=H�,������*>E��kK�")g֪:���_l��x��+���-@[U�������V�8�g7RbV�k�tl2��"xb��>o��?c�f$��N�_�ɟ(x����;E���w���pF߉��d(�y�8�(i��w�_P8���l�y��۟�L�F��	����
u,���ޓpMr���|�Y%�S$௷O3�=�7h��]����kQ�?�-G�l,�a2��I�a:
g�I�-tH�f j���:�O�t���ϒ��zz�/�X N���X	�@����7žc��ύ��v4��~����U���Ͽ���H5���1�\��
�F9n�V۷LA;简��ʡ����]�g���j�����L���w;�5@��F�7A�ޒ���*�q7!�t���EJ-@���T�y�(���j�w�"�`�2&M>�$](�*F*��F��4����M-%ޒdB��9T"��'sk���3��K�D�/�_1H��u��G+ջ����Pw��Dp�>��~0o��ۍ����B�e��u��c� Ơ��ZN�Ǵ�~bLY�<��E�:��4=��PR�:�x#�(�m�0>!��VK��I����'����m��>E�����'�2�x=5���jKg�Ӭ���܁!�����U��<�R�v�٣�U�%TZZgG��Y���&1R,�q6(���]Tv�f\�2i?�(6�J)����q�0#=��/T4d`gy|��H^�P=2;����H��Y(�v�cs��10,VǄ�.~L3h�@�u@A��G���?�}i!v$��Ii|i�~C����Te%|���nD&��'6(xiͣG�ȩ�zv������,������d��lY�2���m��n=�4��UY��R��x�n�>�:��B���t�#���J%UY�)ۃ������<��������\�)>��p�����ҪI�F�g6�ʮ��X�-j.J"8{!к�{���4�؅Ж���2=��zL�����R�7���6�����'��ٿ5h�=ڜE��R�"�k��oo��|�M�A�m,W)��
P���L��m�_��ث9�bX6|1�R�4�/|��,�����#`�X�m6��]]�?z�ƭv1S�<!�V5�I.�z���CCaǗ�r*d�i�s��l����5������S�Ŗ���-n��wVn�)%�&O�,QyΔ�p1p�����0f�Z-3����Q^���x�b�ۋ�%�j1#���r�=�aLtd*��ϢUʹ��i�������oP���?x ��1�K���-��Y���	�k}m53��]�qM�<��7���09�����U���*�#�
��D�b�
�)dAN�x�)�B��&����0A��(m�R_ ��38�h)��n'���B�WM���>Dc�nʗ�m��ٷ����&j�I9�@>~���6�L������#�Wur��ϋ1]q*��^���-�tȂ����!7�kT���.h��¯��M�ǼW_Y��% �*�_Zr�C�R�ew,	A����q��19�Ec��i4JA62�.��K�7D��FN�Y�2�I|XY���e�Rs�n0��.�b�a:����K�H+IMɁ�Q�B�U4�`U�WC
)X�H9hf�6g�`$�c�P�P,|��%���.@�p� ��؍ɾ1���t�_B]Մ1�ȓ* ���ek��,E~�G�3���)Z;r90�Ѡ��g�I�@�e�=IoՃ<�$r�5�dj�ec������� ��K��Ж�2!؃��ɰP����=-;� ��Ɓ��C/Ӈ�]�2�s�L��]�͸�� �l��@n:�~L��J��~���4��]�֢���|'Y+��/+�x۴�.��6�u�`��)�)�r�f$?�/�ܰ����r_��t�2�e���&��8��)U�EDZ������)��B��A5�Ta^�s���8z�Ȃd��-���/Պy���^�h2���bm~�|���:�Ƃ"<2�1����8��9�z��iYqnO��v������N�R��"�2͏�u� Ԛ���g��H�Ϧ�fPъ�	��0��`��V]d���8�u���)�����9�^�Q����~L�I/;�c�m	��NB��7��Xh$9�EÓy�z�kJ�싻0H�e��G}�l�"4��WJ���[���N���D���uӘՎ�Ɋ�͊c��H%�/��ԩcs�1���.!Y���r��?�������>!������z�
�~^H�lV@-�cIj�B%&|T=E۩��m̌&`{q�����Y%_�#��g{(�^��K�-�iS=�%�����P&�`�+r�����ٱ��k*�B�u��
�����e��o�*�g� �P��z |_�*�N�:,d�ޱ�uI�@���7 tY�å�Q��À����E�v����Q1�N}�y-�q��x�=~HD�����6�ɸ�k-�dRuU4QP6T|�WS]�p[" c�M�ˌ�\��}�l����h����T蜈�[�Z�'�p��-��,�ZUP���z�o�������Ϭ��K��_[ ���G�Q�?g�u蒫v�r�׹�)��K���}��:�ا�F˂�����R��GP�&���.���斄��҈S��]�����{�����Z�*m���w1�:Ͽ <��r����x�-3�h5ɬ%<�`c�;�4_Db����g��B�gL"X ��IvN&�9��ΐ��B���!�0{.si�<yS��=�N��~�$�������#�����ę��W�q[�ʿ+	�3��c�9N)��'��nR�5m��|��q[w��4ӗ����{#e��,��g�~SV�e&�$�*�8��au�ki��|׻��D;��]�G��@����)��20���ݭ��w�4��ff5�` G�4�k�t�Q�Y �ϯ��|e����dRH�(ɖ�4�;P�">P�
6�m��ro8m?�9{�I��e�~���ɘqF�X�R|���wǸ�Wh�j4ɶY��_
�@�|�"�0%I!���}d��S�Dr(b�1�>=_��� ;0��ʐ��e솂}Bv���X��p3��f��g鑯Yc�um+4Ss��,���ow����6����=����#h;H8�\XKRF���G������?�A���A}P�H��PZ��R|J�O��)��XG������ve�ѺZ�N�QU`bSk��wf�V����냽����^,�K���]��]A k�SLV3D�p�v
���оn"��>����7�͟R��8@Q�m���j.��BD3�(��:i("|Z��G��ֽL��I�MK`�]��F_[ަJZo�R�/�e(�t��%͞��K��Y�~n5�w�GFD�t>c~����u+.��FW���k�fʽᲃ��!��(*���M��`�.};�	$7O/;�bT@ӵ2p�I8GMv�K��T=uHjC*��̣
;���^P]�����m���1&�FR�'���Dy��gs�V�r�6��SW+#�<�2y�lVxN-,�W`����I�&���kXܝ��L�l�ۃ)-�Ӆ0N|m�{��^��"���Ɏ$���x<,8 �k�;�?�@�i��K���_w����]Y�� 뾐�/�d(��t�/DJ�Kx�7�b�OP5y$�ev6�4i#�T��~�����yj$�
4
+���'�l2j�������LZɤ���_�p�v;
���F{��F�F�FSS�q����K �3Ö	��0� �1񏚑���{]d�D��EU]��S�BĬ�.��<tx������D^#��[#�y�m�������.?�*Ф�/��l�	���;�D���H���E��啇)+�gN��7!����j���@��432ˏ��%c��b�����vv,��ds���`l/a1O-�����c��~/K�
��W�K21�	`HG2)9O������ ���%>���"u3aƝ�BSH�c��>��܉;�v�DŨ/���s1�"�2c��m�ٛ/�0f�R�"����T��á��p�L��2��uh��U��h��چ?Cy�����*��YJ��{EH�;uM����Ig�CZ�?�R@�2�
�>U(9֙"n�#���梉Ԏܟ)���"Oe^9���ۢ4r� �N�{aq>O����"��C̈��e"�)'��m���*AuHTr'�L�~xƂ�4�v��1����т�R�md��Bi*����V�\�Z�jX�y�e��=�m��>��$�|N�/�������θ�� 3՘�g��*�V(��W7u>zA\�]����'c>Ovt�˭���=�;�Z�;g.�SW=I��y}��β�����Cv
Dl>e�dg��H�����覣<u��_ �U�_��i��==�qԤ@�个�2x6�^)*��T���\mX�L��Q�X>s���[��p,��͛M�zH�*��f0C�آ��ﱀ����nHZ*�Ɋ��o��>� \�Kʰ��x
�g�������5-��L�}P-D���3���3�pX��TW�<	)�n=�G�����;O���<���z*k���(	��K3O��1A����^&+y�j�;���[�5�H���}�E�6�Bu�C�Owe�;4Cn���dF�F�& ��Շ!�0;��Ǳ�t�(���3DgGNBA^\�;�NG��13ǧ�?Z��N{⢷��}�n?]rP����i�5aDk(1�M�}�(��*x�M�(,|����y�,�m�P��=r�������th�So��b��E�n�&��(�!�ܱ8�xy��^�*G�S���5� �U�=�G37X��R���6ԅ0Y��w��Q����� ?:F�6��^�NVc�����)����yᙘe)A���U����.~3��_�����:�"�t$qd��7����\1�e��9i��A�,�3tJ4��
)@q}
$�j�Is��߹Su������y�3���VC�CJL�]�Ɨ(�G��Ӌ4����qdt��bl�xG(V�2�@�9]E�v+ �󺺍̎"�l>��4<b��:
 �U3
���D��Up��?w�>������i�!}'4yo�2�2N(����-_ꡣA�|�c�H�A%�J�}�|9z�؀���D*VSdq�z��|�47�t�)�%�̅}� O�_�	���WIr�����)Ǣ��O$���k'V�� :`����uR<F�Y�2���-��"?E ֌����?�yg�Wcd�Z9�� ���E۠��P����hY��3��#-Hc�B�����$H\�� �4�U�L-�H�v�hΝ�˩����6�c=ej�aQ��]��<����z�,^	�f	\����K����^r�� F�Y�vQ�]>��e�^�r#S�8�[P4tw��w
 P��$  �$y���y�e]��Zf��.���[�j�(�C���bD��1��2-c�4}z������H[�>!��Qԡ,���2<�❎c]�=P k�bC���,S�Pf]�F���1�,�^�D2����f�̴�0�̆/ʌ��h�W��Of#��dGؚ��/%𝅝��J|'f���������~Kf�x2<��9B~���i��v*T{���0痌�z����.1C!��I����_�=�^I�:e~�a�Qd[���W��=��[u��G�kU)�+Pt~�����"�|�J����ˢ+z[J|�LnRZy�Vx\�Ɲ������)�Kf�*���F�8��Q:�Rδ94��j�,	�䣽��AS��Ne9�/b�C�h��F{�xyL�g�Mx�$�^�6o&�b����n߶B7�_u�R��W�ז.O���]���R,��K����!�͌���{��{�u�L�eAj����8t9Ф�>�x~\��{�S}��������H�ۚ��{��T��P����clFr����/�t*t��7�Eʴ�k��+�����p���� R���F:@��^�4��d�9�oL�Ђ�Qzva�rI@�Z?�wGz1�6HB�L��� ��L�G$�z�8"�u��8K𴐽	"fH�]���0����F���Ûr���3@<�#����v���`7F�RV"ӿ���.�M&�_���ѳ���2�k?1D~7^��.��ǁf�`m%|�7��7�ap�A���I�h�h���\O��LzG�$q��,���π��2X9(��cn�/���KZU��^�$�9��*��>!�G��7<�j3�]���P��;�  �3WSFX��s��X�/�����8�a���H��=���k��hpՂ��m��z��*erHxգj�ϲ�}���]���!v$�op��
��V�����2��~<+�k��h��7�<)fC)*�q�v�w/�3�聆v .O���������?���w�x�%6l�����ĨM���\Q�Gx)�ۖU��Y�!�y�UX����h����+N����h@��|�|٭J<�,�3�Ce������bZl����lw��jq��.���~�Ͳ�1�?�_
r\цF���kS��;%J����EO���(]�+�BL�\h�jjc}�\#w0\U)_�v	M���u�(�M��f����' �ۥ�iM�]�lSS��t/���,������c:����]�Y�1��$Գ�*}5h�Y�MI
D� �G)#Ald��{�e:�_taR#��a��	��ֲ���6����^Q����zn�ڞY���5w�"�]	+�4e��I��I���@ւ�Lĩ�y�Z�u�
�F�˦c��T#��˞�oX��9E�Y_��:w��c:��`v�����r���9N�"s�STb�&�޹_r����.���bN����
È��a������}�E���xg)Y)µ�aP�Ӎ��Q���Jq�g�M9��R��m���\�gv';�k���*�IR�bo^��7���Oj\��'���B��7@/xY�tΨcILXQ�q��I|�e+=���}8dA��G|��e=@�-]|�lV,��瑩�������q1I k��k0�V����h*�O�=������t6��_7T���~��(����fH,���t�|p���7,���4K��'�
c�������3�8�-�ξ��&O�і�.I��c�p���6M0�Wz{a�����.]��&ٲXm��l���ÑGOF�t^�D��eu�rUOC��ࡼ6�7���M��J`q	��w�B7�@D��&v#�ȴx0c���\���B�Įs�K�C�ԣ%A�3��f���@׌��M�z癒�l����$����t��Q���o,��N.]���v?ߠ�t� �3��7��V�*��c�a�����Egr7�<iVn�-�����HG���"�3���]j�Ŀ5�kx!�ȓ�Q2�'��<�<"�p�w+|���0�lۼ	|���Qr�F�G,^��mm"�âb�厰'L%��Y\ݤy��5Ӽ�;����\+��8o��qz$
�2�,WA�g�"[+W�*C��Hu$���v��>"��_���i'�lR~��bu���`a	�%2+O�K<;��k"��<�u���z��������5���{��ꩬ�-�����'��%V�nk�B��,E����p�C0{���Y���N�W�`�P�g�s�(�K��������UŞ�7MJ[rxmPျ��zN��;��m��$�e_>�/�7��]�v�3�2�Wr�(_�mZ���B�h��K�����s^�ɧٻ�&#E$�>A�ق0�#E�$:Z�������4C�{^���^�$#���] �k��3�ix������m7�k �)I�K*��^@q��� c�6P���'T�_��#��0,R]xM��ų�{5SW���p��x��8\�h&�]���Ьw8�ǿf+W[���[�oX�b+��ӹ�ڮoү�5�_���%~a��p
�*��cu��*�j�7��4ᾃ]���AI�-0JKE��^��+7�q�)�@\��_|;?չ7��8\���{!��iZ��o��s�s�b+�湱��L�
�X�R,��ݻ����T$��m�Q��S-�E�� ��o��'�y&�r����I>�� {�;g�㒜	
Kٵ��hC�VyC[p�*��[_iD�'�l�A'$�:��<ue��K<b}�O�G�p��^�t+�!�n��Y34�T��q�H)�r_j�V�h'K�
��s��{��]$��gÏY�9wwC�9W�$һ�0:s�������s+��:i�6���~H{Y�I���:�o��|~d���������?�M��a���1��u���/���p~L+�{��7ñI�E���-�Ե���1��p���R��xi�G?{�v�1>A�0�"<�S,�Q(G��%�s����h�Be�G.�F�����Uq3/�T���8(��&qp��%:�,ú1k����$	A<\�E�Ka�財�C5~�#J=��|�%������P����5�\�tuz�K�xɈ��q��0}]~aǖo�\�h�lv�,B�؊��ǧ�K�ݴIO��~� �Z{����}��о�ĎO��eᆥ2V�Ia��%�/�x`ȝ݂�tS�1��$���K!����ՠ�c>��]q�Cv�qMG� ŉEJ*����g�#^�m�x腆���3`Y*���(J��P���n����X�2Y]����TG�­�!�s]D:+dߌv��!���y%�if��i���բ�d+��鸞I	��I�$���L��*����)'�v�8ιZ��[)�+�ԴoT�J��ZsM�n�r�r5(� -)�.xi��0�M��A�^؁�<^����B�וMf%9r�>��GF��d�Ig)����$/w��Dn�	�ehG��(EG�a@C�\�m2��ƣW�7E��<DK�w�ĺ��x�/� �
�B�O̶�^>CF��0�[SRz�O:G��R%��h��+m�NX|ޭ�����P��w|�;������O�6��X�+�,Z Y��8s7�

qs_�I{���~�h��7���X(%��2G��I�2w�(�{��3g�UL���r�JO!�g���YG�~]���k�ն$��V���gw��+7�~9��T]��c��(r���}�S�n��W��H�����,�spl�*b���^�o�G�)��Ȥ�^���g�Ƥ���S"��;Р��!Q��Ǔ6dh�G���
��8K��0��m�ʌ���k+x�a�F�h$�.��n���
9nVp=?T��S3�����ꝸ&�|	(2�;��Q�����0q�o�ע�R�G�o�wE�嶻�������`��)y&I���O��@�ǅ�w�=�u'����h0�s's=�߰��d�1
7�o�E��Z�|߬���i��$9vjR9�YJ��:�vMWʌ9c/��!�o� ��qr�|Y���{3��*��\?� }e�
��c�yE���^��z�%��Z
�j�x@vP^��/ι>,9���Cc�PԠ��;��1M�e�Rb4��`����x����ǁ?�1-F#���:LUy�q洞��׺��G�l�	pX��I@쌭�����\����~���Փ��Ci����Fv]'p_�$��mI��Z�`��C���湾Dgm�t-�ºnH�V�=�]g�.�	`öT_��Q���r�ҍ[K�텁���Ϙ�W�=�[�g�3��FZГ�S���01� �HX�8;�>>,� j)KCI�5�#�4����2�P��a,�a�!?*�Y$���{`>��A���7K`47ޫ��\��S��|�c�OF���ߜ��.��j}�&��@�c�"�_a��� �M#&Q�Ç#�
hZ'���y��8�J�|
e�!*��B��Xn]��?"�	.]����eF�	�/�W����+}u���h�^�5��%�]��J��Rr��~�<Q�%�����]��[Z�*e)=ӼB �m"OX/}4a�$�nKO7	��&�/�����(CH=ْ����A��=�k���/�^��w��(i�Do�W���z��KMP��1c3����z��򋝆5o<�8yԹN`m�D��H_�r�nط��Η̭�.|��5|Iją��99���G�����OZ��s
e�k]���`L���Pr�N!\f[�
k��Ó��w8�ei:��%Һy�J�@�Um�� Mb{r���%>����d� ��U�u����h��K`y�Q�b����e�(�Qf��B�uA0��R/�`�p@}��/D���kNkp���Ǐe ����]��ſq��w4`�Ӱ�H+0�F:⸻يa�*� EƉ
qZ��z���6+�p��$o�����0��7�Ѝ|{��\KMo��k\�,���[["W�J��$em{~�[�H
��w���k����y���G��!�ZP��(���+fQґ�j�Ǡ�H��j͒W*����+�BhW�m6��⧒�!q�v灉
�E]
�hZ�3��p+Q�|y[R�f��9�j��E�d��(�v�G*�Bԫ�2]�K)|)����^���!��E~�ߋ	ZfF��:��^n�w���'{9P�Ym�tS�}�@+�̀R��� a����٥�<<ЗWzI��"��AҠپ�*@|Qx@��;���eH�/�����- 8B.%�f���&@߶�
�3ԕ܏"��1��$噮�3[����$��$�;|�7��\��2��O��yc�9օ*=���=�c�\x�p����q���KS �5K�8I�c=�ۼY�{����s���foE�8�����Sr�O�_�Dpa���ĭv�|t��'ɭ �Y�|�X���p��G���c8�e�0"m!Ck��� a^;�	*�oc[BT���~�~)pg3@򮊀����_�>7��V(!2���,Ju��D��?ܫ5�z��2 �Ru!dw����ӝ�i��X�ߧ���B��B��["-������e�	���O�=
�_ՠ̡`�4��-���������$B%�R� ���^�˻Ď�Ћ�������[6��� �ݧRmB� �ih��Zi26�k�aǏ��H��wӌ��VfOѢ ��U��љt���8��uH�mŭɣ���s}��v���7�O��gΔ�W&wa��w-�-i�b�����5\Miꀊ�em�V?nz+lj���%q��yZ~7���b6Z�t|TOFu�wp�Ө�������0��G�a�y£��
��h��w���(��2D�D��g��D��y#�|�-��h%5O����O+û��V�.ieC�D�����f�R\��%�05�(wU6�.�v�T���ՠ��CC�Ĥ}`\=�u����n�Ek��ɓ�#}q*7�áǦ2�'-���!��o�F���:X~^?+�������� dF����]��励��aP��])����T9�a���M�݃Җ��Z�4�����ߜ�Fs%���!)�J��%ڰ��.	G�����Yq�|����@=�m5we�b��	�Yy�	���$yA�2US�2e�����OƗ�ޓS1�!�lǇ�@��U]��;|\�8}J�"\�'�	�w{�_sk���� SL��q���:���ɠú�������T�m����|��_5��A�-���hy�����ʣ������胉�.�V�a���G9@k܂�/�8���X�取��z
�a�����b=ŕ���dd��o{KzB���@;�r#�Nw�Ur�4�o��H���~M��-��d=Ϝu��E�D5-��۰-�;���2��P����P�v�d��S1�O����/JC@߃ ���Z���c�W��'�CT��k���z��Io3�	P��	�;<GyH���V���%���?u��REag5���p ��pC���N쨸�b��1���1�@U=i/=�F.E����J{m_�=�H��G�Y���Ȧ�h��\��G;r�)���N����Њ/8�}@��E��Ӻ�DG[$�sҜp�){�������OdX.7 �|ȔD
�ۗUBN�����C���]�GV�����:����K�@�B�.�W' �[���DP��/d{�T�IXT��:Щ(5��䄎�`P����Ae��`��UEv�-jS|�h��.�@� �W��PF��������0�\�F.�:;k���&�(�=qXq��A�M;D^�Y�	@�\1��7$����X5'8���:����Yn������� Z���C�H�Ы��K�>�=� /�Ǐ7G{+�
��=B�n�+�)#��òk�g]�/^M�����:Z3L��f=�#ʛ��pdo��M��M̗�@I�ȁI�L�4n��S`dk��/�[l/���}�������+�X�0V5r+Y�����V+��]ڤ����C�����ܠ� ��0m�uZ]���#ʣ7�0���(8f�kT+6�'�o'��B��O�=�-�qP��}�'O���.�(z�����+���ϑ(o��7�5m�t�Q&�:Bt��[&�X�����W>g��h->�l�VF��mk$�ժ�Y��4O�״_�����{� *1I%�)�� �t.dleuNa��ٺ�h1�����iФ^���{������=K�1�^ŭ�{�k���<$���i.r�v�k|e���>�_t*�T������b�������_�~�V�?ͭqfڴY(Gj���j=s�G����᮪iŜt�X�tL˴��>v(���S@q�t���՟}Ro��ip#V*��'^�֩Q�v��,����F�6#E���P� �ݳ����.Y7�wO}!xF~#[RM�����z9����Y3�ٸ�9�hO�/�֔��Do��h7��
j��w���ԅ�\$�_a�`#����{�~HK�vUE�d}D~��*����9�,���
V�4\"��[ ��6M�R��?�*�+�V�N��x�4���5\:������y7��{[�fF�P����7���\(�D��{8�����t��M����:���M��g����+��![n�����V*�BƉv�0���f�ͫ����c���#�u�Ӝ`�`�~�"M1X�Om�O)8�V���K�'��&"��1��t�����1 �@$vK�9�V�}�*)��k}L��6�nZ��4#���U��t H,����ySeJ0�ψWv��KY���c�6��v4V�k��ͧd�e�M=�����
�Mv�Ȁ�]�m�c��M��
�Sߠ�ɿ���%�
�[G�<�X�����w�D�$�PJЄ��ҿ�j�����1�/���Am׋�kc�U��Y�V��!z���#<-uBmK�z@�1]�'���HH"�ฦ���me��.2�3�0$��{ �]��QG�C�.Fw�k�U����&�
���O�.ir�ؖ��F�.O�04�Um���Љ3bc���%	/�Ŀ���%2}La؃[s�c^?L2Pd�]Y�x�t+_�mړ����lkYL��.Q(Wv���r�؎/�RK���a�{٬:~�+zk�%��K8�r�RW��j�$�u
l��R�[�m)~|��Ϛ����?;'G�k�xL5%����}@�>J��PP�~�ｃ�fs�X֏�#
ݟ�Ճ�W�$�F��]����8:�$�}���Ţ	�∙��)�I��/��O�gH��q�H�|F�v������u5�'t�_�`�"SS�^�gw�f�j"G�3�~k�Z[��A�$�X��.n��2�Sy!�Icp��`m%i�^�����@��^��a��\~F F�X���:��%o]b�:[M��.(q"����h�o���8H)t%<�6 Mi�5�k���_�B7��m��� R*��+�>E��̬>��P?�2֙i��F8�4C�>�qIˎ����������<��J�۪7<`�(�*�|����\�S��ڎ����8���m���m4}QF~6�W���z�@HXKΐ�%ɰ�G����Q��A�d`P�W8�\�{U����Y>6y	��M��kSէ�"*4s]AY	��Ġ��8����f�1�R�u��$��5�T�Xl[��̐{��?,l���BF�+^(=�O�A�@��${��`R=U�Ms�]g�,"[0�V�H�QѺ�4s��F����ɕ���M*��,�9���j2�Lq��#�!؞��bI�T�e���2�i�Xg)��EN�a!� M��'��K'��G�����d���
�	�H��/�]�Έ?�Rh�۽h��^O��c��V�V�ڎ' w�%�Z�e�q�� =�g��d��;�Q������v��\%��v�d�Ka)7]�i���ls0«�7ؼP��D0�io�/��>�RfR.���̩:�C}b��e����<�7�n�tS�[�ZMm�Ĺ�%�@'��3a��f4N�ys�!b�"آ����!�/���C�$hʤ%�����8��L�
�� 3Z��h�d�5���|πQ�w��J�T�Ǳ�q_�uJa�%Q8���A�q��	5U��4�r`�j�+���:}�HN�^��ڏ�2�r �?�BO�CD�� �;�+�>98q;�40 �X�{pʷ��݌���������5����;�ԝR#�6�5�R��ă!�L���S�C���{��
�t)+J��'0#-�|�ƅ[�:-P��$uyQӴp7�C�z{�X��I��l��숤-���ٜ�M dćz�`�V�Ce������_���	!��{5 �|\�O.��a�7J�|Z��ߡHP��-IDm,)��"it>��ކ���Q[tNM�9�?�������7Z�4ے�^�٠��7��T�ѷv3k|4�jG��:��Z�O&Pߝ�-�ˁ����zc*����?5��6m!aH�w�m�sS���;�*�SP�M�E+�	��*��=��K$t�E|+$��˻":t~x�vO�5��'�d[�N�x�#9c:'�=�Z�Y����5w����(
q��+BB��bEh�.�T�ܐE��oE��n3۝�1�h�&���8����vT{������9��&��(D� �+ܰRNJ��@y���A��^��^줱1N\n�!�0�C�q]�+��1�hv|�yY$R�*��C�T�;�� ��O�xό{��|�Ï��i�.�-�QH~#�cp}H�Sŭ���+1'��63^]�����,�Y�4�!��MѢf�m�W�W+�RU��ܚҷ90k{U$��fD�0����8M�c��ha�M�7%��r��j�����)���@����vr���¨�9��8��(��̳Y��ͳ.���8��N���c�*}��1�D[[���/�Yl��%~��y턵P]a�`�5h=�ֶL!�@D��h�56BA\�4<�_Y)m;z�/�5(��Ĵ�`�����&7�O�S�����I�p���������4%�K�P�9q;��s�v��K4�q6���o㌺m��K|�R^:��A����C��9�)������ة��d=?w�{X^����V�-c�V����o-������Ϥ�ӗ���so����W:�+v��5Z"y�v���3�ڿ��������íoit�bCi�Ro��;�-\%��ι,+H��y�S�����t�jGFD<TE��x��e��ˢ��ݷB#��>�����܁P������@��g/����29��N���f�1�U�E�Z^�5.�ZwI(/�>o���I�lp|�d���� _����ƎlTa[��q����IoQL�0�{�XW���P�I� Ta�$T?f�
['�@#�	_Z�C��x���3_�@17��bZU�ӵ���UF�l�=�`RR>g�����{I�JDF�^�߇_�|_ڹ3���g}I,��S!ȩ�L��L%�=��k�VO�{�m�A���`Mڼ�䮝,�}�
�Ij,Om˘��;�FeqzV�@�T�n�L����ݎ"|��hb�tG� U�v��Éx� .���	�ʔs�)��boX&,�����wbM���.<���*�N�Y�ZmWx�x�92��@>f�/�e ���|O`�0���r�e�����"�е����wϰ����'﹄^FC �Tl��wh �GhW؎�A>M�`P�7L>OG���,�v�lH�S\L]M�U]x�9��/
����A��	��{��v���<B�`)򃡤O��g�ނږ������F��.��uy�Zhܿx���6��9=�� :w�\�Jb���е}���@/�o�ԕ�m篙On���$/�a�`��Lt�﷐��q�@��X��Ym,�Ύ��c��K'O�u�}���ыB=�)�=5�:z=��s���U���_߆�&f�Q��[�G��~�?`�(t��	T����s��c���禇��c@àYm��`x�94K�Q@"i6�&�����A��1 v�$�f����~o�|%�t�߅�W��Rl��i�y?��x&�@�Y�s��ՠ��_��"����K�����ӹ���K����[�U�[�	�P����K4E�_|;�s%��o�"��a��" u�t��4��`ˠ0򐖅��Q�L��Nb7L�q��\NB�L~������V�kHR������Q|&{
��c+謶u�p�-3CY��N[M�h�W�Z~#a�(�[-	o�������"d����M4���7� ���]P���5rY�"�C	�A<��0���^�R��n����ђ��y㬋�*x-��[�> þ�XI9�6��H���[)Jp>��\`�FZR�� X�_y�%�6��Z�/�r��-�,���=gŊ�g��4��kw���'��߼��{�P���S���[B�28ό^�9_�EO���4�O���]5��R=�SZ&����!SRv0�&�w���F�e�y�_�6H|��B��Y,��6�j�at[O��e#O���?:g*�4������]fС59�ML��FV*�p�J���,G%0���,ij��V�q����rm��,<K ���3�B^Z�"΄9�E��Z��T_� �p�\��gC���^�N���+�_4�O�٘A�[[�J�ORÊ6�?���������g����4�T� 4;�|`ͳ�s�������uǡ=c�it�e=�1�
p��xٕ=���]��ja�:'�^�A�Y�.��6v�<a|�����;��O�Ѹ���'c���E$�?X������N�Xr;�����Ō�[�@X���0�k=�M�/�'�<�l��[������R�s��q�,%9��b�|�ڏ�^<w�5m �;���X��|�a�d(�U�<1O�v4�����(�!���+=��D��"Pe���zW4�" o�*Z���"�������>(�Qt���$��&Gcϣ��
�s������H���9��x�����{�;2���1~d{��ğ��d�̠h]����(m�p�t���A,Ё����L�6��˧�������vL��J���4��,Qƫ����~>�~�!����c���Fܮ2<V�ItDZd�AH�w%(���FD���B�R�a���gĝ�;.T�κp�b����h�"U�ox������F�l2T�T�)�F�WaF0K�I���B���wT�X��*e��*�w������4��3��� �y|i�l�>�Aq=�jٚ@%�6�lL/�@��R�̢�����k��S�"?q�ݞ��
F�Μ`��glS%�!usO�@.�^��ש�&������W*k�e���C;���QU^QC}�Ħ�r�ULJ��Y��ְ��}������h-	�v����Q#b��
Ьc�����̀厛4�`!�hJs&z�-�s'i�����R*�an4�����~�t42q]��a�G)6~�I�5^Z\�q=�Mk�I3���節fSD{��*��1ktE�Ǜ��g��-�� y�>��ll�E
��zV�ȟU7���d�MY���xeW�2�z!��|)�%�HM ��Я9�>�"����#+8h=�V�֤��S�Tjj'�(�|���۬\�E��(k��+�f���va�s��zv�P"[�X���F��-�$X�9�B���8� s����3���5%/��f��(�6�h�f6��C����n#�q�?e?��(3�d"�`�A/-��_���x�\�	�J<kom����P|\���Ao6����,����n��\$]�9S4׸/�!�4�դ�(6����g�[L��^�jz&=��i��>Xi�e����RZ]!�2�jB�oi�t=��u��R��8��O@�t�f��N3���	+��rk�`�<Q��D�L).���K4zK	�d���%��e!���ق��Snˆ�`����q�a*'�E��1na꥙ǅ{ֹ�L���=7�ΎjO#����7�^�;0b���S��L��_�r[�1���l�V2aŦ�|�1��B�Q�����jw{���r�����
zc��k�KkZ����ڼ���G'g�q�n��kϜH9����h�K��M�T�.����멅�b�0��G�7:ɳ�w>�M�h<Gr�,
���}�FE�s�e+�o9�YRu��m�������{'k}��:H؎gv��Ԝӗq$x���O���ʧ �r�I.SfV]��
�������f�4�%�SY~���v4p֦�Q$�N�;]�
���(=��;B)�v!4��r��bOqՕ���z���k�O���~c���b��&:���h|�*#�^����n��dO�nx�\��*�Ig���2�F�fZ���Z� *E�QI������+p��/n�2� �/��"-�eW-�]�u�[C	[��R���O�+�><������{�i��T�h
����H���JbsB<���f=� �c/�%(O���;Jm.݂-:�d�D����X��?"�iܪĪ��&1���~����4��BC@h���w��P��AP��ؕQSm'�]+*`U`�+�J�؛��=<����-X��c�K,|������U�3�lI랉�
H=�Z3���s�"�z%۰�S�|��A��G�z�J�&]������TK �'Ec�/i>�1�*��9�4֦lJ�4�4�n90dE��GG����I�?�/����k����_=Ҏ)��9�tP� z�f�{�ߓ��*�8J�Wj��H�\��$
z� ��f[fb��Ʀ���u���fA�7�T�I��c)<��°��m�u�~cR{��[�ۡ*�����6�r��p��IW�l&���.��Os*�p8O��"�z�|^����I)��I-9�J��'�uA�'E�6��H�����l��te�J��ٰ�I��p&u%~�4&� ���5�h�bg�0�?�_h��b�Y��s�cO)U��E'�ץ�#y��=�ʠ����LR'oIU�s��9ˍ��yN+c��ޛ��R��f	n�����?&?յ7T�]]�^C U�eWg" �_����66�o� J��L'��S�	O���`�v~�$c�f�3��*}�#��n�G�!p7\��d}�S�ښtq} ���Pg�cW$���9E�S����v�)�$R��`{�֌n�"�34pm�0�`��5��a���/8�*����ܶEeSv��+�c�oe}f����߫���:G�t�?�Pj��3�nh:��#K�t�7��Vqs����s9�r���)d\6ߒ[���~l�V��R�jПhj��N���/�(�[���|��Tsg��Ti��K��kЬ�ARuK�9ho�����?b=+2��B��!�Z�i�sDĔE4�q�����S����-���N��c�r<���4D����~�Z��^o�����k6�5	,�~oo+I���5�a��ij�q"�A[!�P����F`~��+��8�R��{��Bf�Ĺ�
��SH��\!��o�Y ��.�QS��@TV�_f�v�P͏^��<-+�&
Q�,�KX|ʅ�X��f�1�ʙ3TKάϠ��t�H�L��"Rx� n�����M
��y�O�������(����m"[�B�7�b �����aO��\�B�*MLm#議�SR��=�Z�������x͑��S)��P&,�D��E��0��zXg+Ѥ��I���O<^**�5�Q#��[#h�@ɧgol��������K5ޑ�0��tEN-���>��@�%��Y�{�K��?����cY�19P��kU���'��mc�β�A)_->�@��s������ ��� �zO�vn\*�K6s���%d	gs��F�Q*�E�a����aMC��:+��� �����s��ptM�*ǒ���u�>v�>�>�<a�߮�J��6]�N���1D�j�[p�ғ�"D�	c��F�ϐ]�h�vݲ\�/U���E�.����ڒ���m�����]�%t��2�믗�(�437x�Ńx1�E<۬k����wd�1�3�f�D|N�w2�	�RS�i��C,�k�V�w������$O�@�/b91
2M%��͒5SCX��mŨ��@��=�@-�y���]�L�$� �����;�T����V�7��,�� �q���	c2�Ȧ��F&R��Yd�\1B���쮋Ø[T��>,�N[�w��m{�y���>����(.��{6�A����8R�l��|�t��y.R�+l�Ә����T�k|��&�iP)�2-'I��o�юhS�Z�8[��\��P)��ѼẲ�<�R�6N�~p��=�ii4��a~	�5���_�u
`9�sy�yZ��'|0���'9����ܒ؎�R�L���Ċ��/;����Ǵ�`�F�T0z;w�UbK�R�������i�?-�?��Ώ���8'�4X�Ermq���S3���3�� ��I�GM���3�22��҄"l� vE���0V��E�tN���\���׼ڏ�m#"sV�������c˅� ��$�a_k����`��7p�<�m�%	���v�fV�#��hOo��ly{�M={X#���-|��9@���	r��!/,�ӵG��Y�|�گ�'�N��}���{�0�����U:C���_���h2
�5�#��C�߃7����@,�J�3�)�+
7}V�V���Q�p��cOt��)�b_��������joM�$���2/v�ϑ���I�0`���8e����c�:��ne�>Z�B��I{r=����*>Ѯ�c��R�᥾�|�ڹ.jRQ��pY=�j
�K��Jp�u�Y!Ik���{M��ZfYP�f>�������f3��lg^,?sI�xQʝ� ����L��x45�L�d���yj3o:- ;߮���KM&8���2y���m�D�}8c�vMk@����ED󬻙T��0Ҋ��=V�Ʉm����^0'�X̱�rA�a���ȂE���Ӈ����o$o�����#�U�w,�'���k��z"8�Xt�<1�E@+��=�� �Z;��7l8���y��
"W{D�z
9���`�,���s��c;�S6zѲ�+ oh�9N�ӻl�ޠ#�#=}��!��L�Ƶ�����*�B�_�)
�Z�z5ₑ[��LwY�T;t���l^��X�뭠jW1��J,�!����V��-Ӕѹ�}$��[��H��˰���śz2pr%�.P3����GQ���²D����s��2e�����~�	�A;SEqTě��T�/��ه�4�[CF�#Z�ߴm��q�������dM�7�@���v)�fXI�~`�F�79�y'_��d_��|l���W'n)�)j[�4�#|e&h��}�?�,��A�P�;�
�L)+���ә�G`}.	�Ҽ�B���'ڻ� eIF)�v�x�V�3\�]�@�K����pqp��O���@���xRG�*ej;A�	2EyM��:D������l5�}�M�~���m��HS-��ϋFX�6S���'~���_qN>��~ �v���P��kuq3�V%��e��{�y��5��?d�� ��S+�����=x��e�����S��{���e�DyW+���|Yci�&�]���Ľ��,Ӥ�7s�������{����*����'>�u�NV�A�Z���q��J&C�PQ����c�-����ԍ��l���|!RNe�~��}�0�3���z2c�5�>���������]�.��=j��w�+�e�=lS̢�kKP4��v5�4�G�!�9���U�!`�`|9ɱ$󚽼OO�e�K<��Y1�#a�����g��wB@��t?���h�S�.Yf#V�3�}&�Ϝ[A���!ļK�`6�g�\b��%و-��o�y�cs��-y����,<Axo��m,���. �.��Ĳ9�7���XTb��d,�A�	�vH�r��m1��&��V��ŀn��#�z��ڒ�?��kH�4z��P�8@�V$���?�:4��m�5�ф���6��m☫C�z<h?����%��$,φu<i�X�����{q�:�6n���'��E�+�d~��'�'��}��"0=F� ���ri[a:"�@�agv�E�t�ݏΉ��:�Hm�<;qm!��P���2[�+#�p�	��~���'�5x���0��qXw��C��RJ��|=�~�7�
x�Sl��Og��í�p��D�m	B��<�����Ή�ٴ
�.)�L�8ذ�#t�c�6��]�UT	F�袻	X����g���q�O!�5�G&���W�+Po�ǅiL��d���r�G)w#p�O�uB�uh����B1̜�-�5�@29��G����[��k,΂An�Q���E\�@�e�s�_5�&Rf�l�d��<�ZO��:���b���a��أI�rvi�5�+"�s��~���@�U[,i`^Z��E�=��5 ��0$v��vTQ�n�v���SJmf���J�q$f�0::�'�2��7&�O�G��h�T��~�0��&�W_%����9V�4�ˢ��Ӻ�Q͗����`h��d1��?�C����B!VF�Z1� R�Z�� ��=%����zaiթ�dá34g�'�+` ��D~� �>��V�-������~댵�jU���CI�GƣfG�J�k���!�(l��.�D^F���D.�索>ǣ��YoAr�����4�1���܎�t=Ԍoc*̃wUWĲn�RQ?*T���an�כ����S�����ӑ2�=�E�����VinY�V+Ӄ�][#2r}��/��f&�9V�@?g�ps�%m�p{8��	�����}��N����ӃXo�xέ�wm�*��p���U-
G�����^QR���;�_����l��S؜�l��?�����AQ&��e��|��i���1c6O:��xxЦ~븈"8ANb4��P�f�&B�	�'~qGm� �X��6M�]����B)�(��_	����^tǎn���J�e�ӿ5e\3�c�NR�B�k�'&;@�"-����ϝ��R�Wk�@"3948�=w��ې��֭.A��J��<��2ͦ�����Eɂ��00}�
ީ^������ݮ��B�p���9�t���ȞE	����F������Ij�p�E/�&��<+K���LY��J+|K���]h9m�ܣVF�qe�Z�q�h�q���h�b���5*�g��L��*DoI��p��c�7fE;��I7�
��z�q�cБL9��r���7��>w������Ŏ>	B;H�\T�=v��R�p��0J`�į(�7�ܛr�0�-r��	T;�e��Z�n>�Ye�Br��:����!L���BW[����d)qu��@�篔��#��l2]=�5w:�B>kU%��g�u�h���U:��הT$M
��)�(A���Km[-39{0��2�N�I�d�*K?��o1�R\<%�)�ş8G����ſޖ�3�:pB��]� 7����r[R����|�%�,�h噔=WQ��(������Z֫����ĺ���E���m��,�����N]�/e�*r�J��e3��U����pNK�jz7����aWx�$T�̓��V$�(�	V�C5�|���,Y�e=�	l��K��_��tu�B:����Ev�6�@!�7iJ��s��Q!m��=�Om�,�$�,�<g$Z��n��w��������.��}"sc<i�L�g��r��He�KW�e���D&P^3��1����+�BCp����X�+X!�\5&*2}e��9��y�+RM7n����ē2�SmW
��`�xK����=���Ö�r" %�o�>4��)���U�\ ނ�l�s��[P��Tt��)_�DV��ϡ�mo�ZBp�)O����L:�ߏ��Z�Ⱦ���[^�U���Q�PЁ����"&��P.�\_
��u��^�`��HU����E�VJ�M�'�y?e<��D��bH��Yܕۅ��)�a�hp�V�"X��Hr�#��,�6ԝ���C�z���EE��C/�=._��*�.�VI�JL�$iR6�r"�Q�~DT�0�L�/8[J�����6�&�@�磟Dǂ]r�2d�u���-��g Oʹ��L�r�P  FH��7�@���BC�C�Hj|Rj��B�Խ��;Cd7Qa�F2l �1�`�&�F�(f^R�}SrA�$
�-vM�vW�� i��Ƀ!OL��i
��EK�"�z��I�W�U�K˰���FɌ2L�2�Y,n����0��g2Ϭ�va�e4��`9� }�����W����9��ַ�AD��R�P�o�.��ƫ�Md��|���`���,�g�;d��v��C��M�#�����ƖY�\�ܣ}-"����eH��R�e+���w�����u��Q,��XqM�a���ΐ��-Bb3��@���$���-<���@@Z|CAE2���'f-|z�I��0�2����̈O�,�Y�)E8��`c6�*	���2*�fER���-Gk]���G�v��j��@Y�e�F�]�㴶%k��H#o�B�8 ��x��R|*2?8�2IL��^�4�f��_�	�8��7F	�K!41U� �n6�-@Z�k��<��1��p�Yl-��t}N������������ ��y |&k۸�a���w�~+�,2��v�妊C�����N���T�ߜ���)D_�5�ډtr�H�~ $����#�u��Ot�2�Ǌ�4�	$b0<��K�:���u9��5Hy��;��0�D���ӭ b��+���cx����ϑ���|�:�m̻�9�~Z��̙>�I�e��+��=�
��t��͊����Hl�2>t킏����ok�A��[)�>)jU��񊆍�-���e�%��*�B��H�/' �92�C}�{O6n��.*�s�H
,���q�ɼ�l��|�2�т��I�[�'�;�bǬ+̳��a�!�hhlR���\.+��L4�쥽+m�W����(��~��Q�%Y�� Q��W]qz"�|��.-yY޺��/dA�%1�u�tD��P"=A��>��q�&�<U���pHJg+���|�E��\���[�N�="���,~�G���̒�0�6E�Ql���/TJ~�%�;5Έ�PF��<;��o���Vk}d��B\6�PJ��y�`d6��
r� 9�$���:8ҕ0��n���?��/$� ��"7�(� ֵӚ�&���?�X
�n<�JL_g�f8���veo ����8y������e��)���^3��?:@���{k�/$˥�K�_�D2:a~,� ���_;KJ����q��+\` �
퇈���},��3ڥ�N��Ɗ�TEԉ���	���2�k��f�}�4��HY?kO`+,�M���[���2fd'3T:��!f�i��)xC���h�ڨ��bLR�d�ہ$o��
�b��`b�H�g]|��Q�jK�}���ߛmɼ��B�-����s���X�.��8�u�'��Y1K��P9�[z�	�y�Rv[��-�"{�бL�������Q�U���|�,m��i�O�8�L/#���L*�X_��d!sۚ���{��q����\*ԇ�ϙfv�I�s�&	Ը���R�90��n(eS��p���zC}�O	�M�n�-<-�%|��� [e[��,m@�Z��@Qvq4-���3])u|�18j�n�h"qOD��`R(@"��H��&����qX���[��5��|N��p��.�_1���c<E�	�nv����@<���M7��i�����!,�������V�$H�"2Fr��!���*�'��\ i3@�K΁����_?C�J6|�8���2*��3�ZR�!N�� ���C���sɟ���©�u�R��٭�7��#�j���%8��8Xc�ژ�dWdE��t4o���km�
��|��B����/�NW��H396�[���T��kϏ<�JO��'.+����Ǖ�T�3�b-t�$�Mۗ��g�f��ŐMp�A�$@�Ń?W�y& �/$�*��K)0���_yZA��_#�Q�a�
�˒N�b$��Sn^�5���~-�y����J���MF�k�6�������V��9��-���-� ndP���_/�_��-4�p�q:"g�K<r���H����������K�g�������~Jhs{�M4D�3𹾠����̶	71�L�AcEWi����%�=�߭S����� �㍍��
��6�����K���˩�eoR����!�5g`[��x:`�ui��ms�H����{Sz�o��'.�3����͵@���r��E*��ڶ;x��wR;��;�ֶ/Dy'I�ϭgX�N�G<h{0N���X�����*;D34Z��I�>�S�u���
���$��Y���i��v�`id�)�;8�њh���)�x�>��D{���̗��WI�io��Uʒs�h`?��@U�mz���� ���%�o����k�����f��U8Ь3���wK()����/т&�!> 8q�d�~e��f��^�Z��~�Yv�s
�+k1�&2�����z�6���	qBn�����8SD�|�a�ڃ���6_V(j��(��ѫ
,=K�*s7g��=�4�G~������Gu:��(��Z@���Sb8�1P'���}��{"�H�B��*���S��Ia
���(�`)��Ab�2��`�4��Ӑe١������*��x5�Z�����\.ĝ���дު� %�_x^P`a��̓ ��L?]:ȏ��T���a�2�x�1I(�
�F�����h���X�yB�]!p�3Z���7�Kb���+Q���A���C����Tj)/.�VN\��o3��\�P�������O�~vzO+�����q� x�X�̮��ڻ�Z�\�f�x����1�RE���}8ΉBn�+����k9g���ϕF{�z�N��:�l ��c��ka��۲�rMG��O>UKJ�J�qͯ�����܋n+k��5L��&(�2���s����ڿ�a�<~E}�u�GJ��އ���rK�1W$�����j�z�pt�bͭO�r0���e^��������,4Y���'(T>�/ݰ�r��G�ߋ�>+߈w�m�]�>̈������p��$p���g�[��}�����<3��k�8x��N���lA:��d�5WO[S��9G�"F^�Hy�a�Һ(�/�`LH�M�����<&���3aRw�A�ЂE�eޭ/r�G9�5��Mǀ���S��Z,�%������"P��Ru,�j	%Ԅ��z�K;���<�T�Tl���0�,�nVQo��>/r.u𫆹8��4��]�gS���?]��幚g2T��}a�����V��؆���W{mܙ�qRP��	8-z�Z��]���oe5b��p<�)�b:H�7�Ɍ[�	v�S���=Y6���c��2�	 $�d{?����sPi���ȋ�br�R�.e��x�/`��U��Ǽ�󌈕��"�]�ׂ�RV��^�����#�?{��Qh��Z�����'���d�R�Z�U�J`��NɸX��4z5�ɓ�RnQ����������!}n�r9��ם��y�B9�����~����GK�pƥ�:�`�u~UEdp�l|I�^딹�9Z�V�3�BϾ*F�s��/"���P�;���$:���X�i�a�y\B�h�N�ݘkK4�R�i��ߩ3�aE�-K�	[��aw�{=�-�d8Xsk�[��^b��iF��9o���t��<��������f�ܱO �{X���b�w�����7k�,�7����2�ٲؾ��\R�����/͉H�n�މ����Bx��ڋsQ�&�A⼐c��!Q�[��3g>9�<�-p�5��/��T5�#�>]۽ȵ�V��w�:�Mp�?�l��%�^/3MԦ�k�}�@�vIí�����f=�55�ip��Ί�p�j�V�d����e�lsz"��@�~хe�����E��4���S�L��?��m����Čs�����9GJM���oK(~iמ��mО���=HD�b�v���4ȡOy��#��*��2���=�:���;xeҷ6xh[�,�4�~��?��^7����/P0Y��}�\?٢��1CtP���[��,�I�h�O/�:h�R�ջ:��Az4��m��r��-I4Ř�f���N!�q4�DDy�Qަ�(KC>9�B��\���ʿ�r���!�����1Ҡ}�Eg�%��[����@��&�hǀ~��ն�<�N`�^�ŏ����o  ��<�ut�mة��8������%�it@��a$`f6H��|�y��#T�1��f9���vCJ|Xh�᫤%�����!Ƅ�m�ӛD.y�И�H/�U��2^%ɍ����|�N�����)~I(��w޼M� �����Ԭ�{5�����-�>�����HS��~$�e���/��\�N�A �ҡY8g��w��|�� v�я��6ݤ���Pѭ)���/���ߧ��ݏ�8�)mD�B"�J�����@B����C�����-���Wh&'۠���ǲtQ�4<������� �YS>툭�`�_E��u�H�K�?���I�<��N�
��/r�{w�6d�������hl}����p��Y:S�1>�kI�>=w��2�Ĕ�~�?_^+�>�<�:���u�4�s����Pn��l���P��1��e�"������O��S2�p͉����T�|�8�����g�2����J�w�&��\j虦�9A�"�Z�G�7Y��y9=���_1��8����%����{n�X-��0����h��o�S}�`1�:ނnV�`W���ņN5��Y2���o��_(p&PDu0�����T��i�83���� )���.V�6>��1����T�����@�&L��Ei�h\���9�	�O��y��
�>R?���� ߬����|�R���GA�q�`{)�)��"D����w�4�US+; j�|�o��S�l{�3��n��Ee�g/gH8�1kg�K��B���)�4�C�ǲڠ�To�ޯ�;-O�4I�+��fy��/�=��T����]�	I�ӣL�d9�X�$$�#���NՎ��(<�P-�!�މ����p7򞷯��].돈�r�/XZ�)��$�}껖��.	�_L(_YGQ��N�-���ҹ4����9#�rNA?c|�|db��~�n�Ԇ��_���Z�#����a&�~7� E�g/���� ��8"d����]H	s-+\F��c±A��u2�@�<�J�y��łF�$�h������Q��*����gE�N���Ǩf��h��ŗ�ET�#ͧR�N��!pJB���͑釩N��B�=�wr�I��?;����o�i��t�c9:>~�y���I�x�S7��Dw1Ɣ(�@;��G���"�!�%����=G4\�S�+�!OV~�F5�O?O�C�-�!���
�>L�1�����+w\�JwO�-���-h4e"�}.+��1$t��1<ح迱_�&��^��Z�2,�Я7׀�@�rk�^Tf��4�$��g�ev�G=#��S��O����*#���ξ��(/�\s��c�Z.y�bv��,��(t&Y���$���O7x:r^����\�����`��`58f���6-�S�-��{t�EY�=Sw����ø���c���-��K���Iם��a��F�� ӆ��OA��0Y<^�'ǩ���L����'��d�أ��)%��!�.cD���r��"-���P�m��)6I8/��S��7�s��.6_�|�T��eo�g����&/n7Gf�t������H��F�N(>�9��v�n#Q���CS!���|��8��ˀ|�QN�u��	������	�%�)�x�1v�)�m�Rs��C$Kx�;��X�^|8�D!���:�U��b����z�j��%�`!�oˢY�?]7�b����&9�a�DR�Xt���B��w��P����)����_�Cё3��q3���-�[���"7�o�r�'n�JY�2�+�5l�sr-�4�ka���֠���\䎻�r�*4guOc(�~�kY
{�3����.�3�{�@�:�"g�!U���݇��1�����B�7_������AO�Dv��Ll�ؙ/�D�#9�IK������kg�6���--�@����^�h�zU{6C�����[+�4 1�`���Gü@Ќ�l٪�4�e��#1�<Xhv6 6��p�G�(k���x�)�0`%��T 1��i:�w/AuL�{���35YAU�����|���+�Wv;r"6D����=shkY��:Bt�ޣ���c�Ϝ`�"ք5{����VX����%?�����Q�o�2f@b*���׷���	�2��(�vD>N�rE�����w����~�':�I�e�$�YZY璀�j/��i0��05���y�~���+$(�V֒��6@���wU]�"��ri��7����O���zY�u1��I����X��89�T�!�Kߟ7�F˘Rs'A)Zؾd9����k%��8�HwyMn���vӬ8O�Z���GĻ2=��AAU5�zah�D��@ ����m�Uu�V��H�4|��"�4Q����H��zM}+{�F��p$w�v(��R�Ę��?"�7Dn��ҧ���:y��9���et��*	0��؟}���Sn_�zo^�u�@��k�N\xkc*;9Q�D�7��Jq��v����SX0���.BNq)�QQZ��Ƀ���33����ZO`&o�?��-W��E�]&�tS(�����6�h.����
]����(l�SaYN��0+�5���/T�֎,��;�5}�(ATe�2k�Cc>��]J1xW�V�l���̿+ՠ(���'�.fsͼ���MS�����Q��n����$Nͼ�����Ϙ�~����h��R���mZ�kzMN���.;�?]jj�\�JM�)I)�J)Й�J>�n��:�`��s��&ދ�������c�A�RP���3���F���4)8�ش�Vڗ��(�$�����}����&#�H�;%9nf�Bt�����a�scó�����@���(���96�Ϗ��"H���㼰�^iI�������͎��	O�ǍHO�������s�;�A��`_Ȳl"*��;��"�q��ǜ1����t�$����P#�p@�vl
UP�&�(Hk,
K�߅cV�ы��Է���� '6d�`Å��=F	"�@�y��^�gǵ���N�\7�zz�l��߻�&o��B����y�c"dL��_n��rdP��qpC��:��>����3���'d7���ʔmN�PJrSk�4kA�[tW�4EDW�����J8^��bY+Eߋ �?��*XR)�>�J�u���g5r���Iމ����e<ɠ����;���������L�����[h�&ÚjCڧ����£�!F�x��Y��-򦓦"���#3���xֲ�O��ٴ:a�d�`L����Ke/�Nw�������O��޲�3]d��;���\o����֛���{D����Up�����dx3���7a^_[
�@�)�u�,�S��-�ɼ���6hD���"�
�Oz��ъ4���::=.���q��-�&��x�* y����@��~�2�"��f��^v	�	��m��(F���S�3=�Y�b7uxYu�M8�3΂&��e9*�BY�%�jA��>�H�Fbݹ�33�,e_	yA�!�7���m+e����}�c�d,hC9��w {	����e�H�[���`���I(*�u��
��c�Ss8I�����ta���R�M�y^.�Q���}%�jw�^�K��#T�ID�}���`m���(�;�nͽsL:��{BK��ӥs�V�]l<��$\�� B�KK���S�4���(�C�C�����1^�o �9�����O�:�?��E��S�/H����Ďv��U`�+�Mp���z���8�^J0��/�'2�Qk��~��u�v�\ּK��H�����e�DR=��T]���/�Uү34=�ɋ�b*,I[
x�#��xBHEw�1����e&�|�N�#}rI��-�:l��W��Å�3��S{���PӃ��=�U;H�1��Zd�.c��J�*RC��`x�Qhpc�~~�����巻Y�����[N7�~�<Bb�9�tx��~���WpZ�w�;tF[CXV�D�?9:�/R���)����&p�N��eCN/�����g@���{HA�~�e�},�yq�V�}<;E�;nL����̣�}��g����(yU\��/���p�\M9���A����Ȑ��4X��j-H�>T"�_����n�r��U�U]���ޖ��.�v�Q2u�@�����?z���qv�N=*a�Xo���t����-�Nɕ�M8��f'�#�H�bǐAzk&߫]�Q�HQ��xP����5Cc�~ww���rX'���~ݹ��$ɑ�ގ�eE������E�o�?������pMJ|�BR�#O ��Sף^Cx�-�4S�+�w�ߴ�[G�2ٌ��RZ����䃛曳�=��U�[}���s��F<�D�i;_Y��'����u�͸
�N��/Og�_�c�˕�f�"���H���&��,n`�A�U�#e��W �"̇R�F��&t���ƕMȀ��@,��n�'����}.ݱ��<�̉���=�B9��_�FJ��\��T�ֽ)H!�k*��2����M�\��&�p��A�zjT�b�H8�V�0�a��#g��T6ؘ�܋�u-N�i�O����R��M�\tFc%�盝.|`1��3�p�g�V�d�?w�ü'��5ik� �nV�S���](�'f�������7L����`�����C��M�ۭ�>��>�����;���hsJ�x�,L�n
]�k�\�ۙ��;�;�	��*Hg�u}w+=�u����R�ITM�\���<��T��;k��E�.�%S
���s)�lJ0���FRG��g^ɝ<�S�Prf �J�Of*�z�.s,����i����L+5�d�rhFw��@	��U�o�7ʜ?�n��\[��ҕ���j�2�T~3����d=��)a,�z۰\9O����q�rG�B��Mux�&-����6CCf�'�@�Q���;��1n��<ѝ��F����q�6M��6�7U�X�^0�;ṏ�/ѷ�C~�`�Ht��!~�4�A
@�X�;!��ʕ�>��|u[k�b5���h�jq�����DTY`��I�s~��7�q)`*儇�`��=Wv�S�\e�2��19��O�Q�`���p�"���Y�Qj�9`����9��a�Q@��K2G�����8�����<����ڭ�DN��� �_�Da�f��� T�J����|p-!Z���4�)pC�R�Dt>;>���,'P9��p���g����I�o
�M�e>�;Ļ���o�0fv�p����{*��V��G���� �Zp���sЬ���H�.���5�P��s�'q_H(��v�`��C�q/M�� �$�AŽz�D��z,Ѡ�ޒz�Ņ�?G���i��fiD%�2��{�rՑ�5%p���c�E���z����	��:��H�t>��1�����#������1�q�O�>~-+T�k�Y?�|=���_�C�m��D �����O��P�_ջt����+�����k��7cR'�a	S�|�l�3�u�ZFn�����v�B'4�|�ĳ(�,Aa��*��)��"�̱��MD����Hq��J�I�cVV�*8n���4o&�L��s��$���۫�#UJ��-��[�j1��O��b��f��<U���R�����w-|Ez��`�RRܡ�dX���j�&�*��Ѹ���B��b3��Ÿ����<p��#+S��j\ޓ-,tY��<	�8���=����&j���Z�y	'�V��+���*K�S&Fg�,@i��Ox�{�`Er�V���e�2���c�L���DX��p�SH9@b�3��g?N��7Pq�RX����VS>3�᪡�ǈb�Q�2��[��p�)��i��dq.4.6�P��#�יO
V�in�}	�����25�����=k^-���Q�[x��k�p7�N��$�H�F:�T��f	�[�E���$9�۠o�g��Yk����-����LP�57q�?�(���[�%�p���HZbB���������,��'��nHg��Gh�BF�������2(Ң3�pg�T�sS7����M^���L � � �%���x ����HV�x�ַ�� [�,,��,���f��Q[!�z�b� �
W�9!�E}��4�W_����!��(v���:	>�:��n����!��#��gs�+�����M�}h#��'&�c�R�{�X/b��X����y�5!�w�[�G���T�֛b���
��7_��j:����I�q�L��)))r�i�p�%�f�����
����0V�:i���K�;mv�]�"���Q��4T��D���0i�:�,�7�w�A�խs8���xj�����1��_U�5�I;��?�B�}]�S��#y�h����t�w>��X�*t{QrI:��z?z�b�:�	|��Z`I�9&�\-�18|G�91�u?�]��m% ����%����O~��.��O�wm��\�h����qlA,U�!�^����s���I�;��:�t�xҶP)L �s��x��$�"��ZO�%_�ᗷ�s%~C��~X�S��{�ݺDEs̟��-�^���,�I|��jQu#3t�2H5��I�O���=�6`q�W��M;ϑ�J�k�� rt�7���/��:a���`c-)sHӎ`2fn~fZ��*&zA=���/f܈N�4�Vܲ�j|�-Tz�g�8��r���0�֞�|�b�E7;�����dl�Ø.�Qr~��W�ae�C��v	;(��S>���(�[�X���0t�{<���Ax&�m��1�!����Օ�����G��x
�7?�����b<耏P�R���/��j�aj��������^~�9�l�$��@R4�u���N�ټ�c��G�#�\gt�	=�q:��v�]��m�w������G)e����:vӏ�N������KX>0��2yM�<]7�����/`p8G�Ѱ��T��W;\*��R�B��*���h�az�����9;;�u'�@��� �ψo���P/wf��*E���Lu�֓y~=�D)?&�J�= v�C�L����ȗ�?��U��9�}��,$!d9Fj�ځqz9(=����g��ϓo��)�����`X���\I���-�DuT;�W9�]�������e�ֵu���G��	��XYĖ!7�3g��Zl��멁�v�"��/�md��S����b��np�Y��u��z��(��.Z5�I��SZ d�1���ZS!"4��_�3�|��Yl�Rnd8k��12�ý�u^r|kD����7uڪ���;�;�J����Ay�퇢��j���F��Wo��O�I�<�8i�w�&1hb�$��956��� �'�6��&ͬ��98�=�����}Uռ�\s��7��72Ht���Z�-���[��F	G5��T�����N�!c�IB	g��B"�y�qO��O����"��rZ֣���W��<����Bm	��3I�kw�w��QU&KZ��\��zL��}�>�T*����O���0���cn�_����[�תY��z%��?[n�~�y'��>���KMj9JN^.�B����s[�⢈3��R�d������E���W��L=-S=C��p���>�xD[8N4�K[����B拦N-4'�0ZS&���v���J���7K��B���������
����t0 �%WId���a���?�#/����p�G�H=ij�TIk�O���j���0�����}(�g��_��H.�pX�C��G#�E�f�㥑�~��nܲ��)��:&=�����y�k����2��~�[42"�`�&�\��;�� ��ި�8Hl�^��>� !�֩�U�4��K�xSz,�YP/a���5�N��
67:�]4��+F��͑�%� �O�Q1��d_w��������l�ܩ9���Ws�)�۱-r�hgU��2t�&\�n���՜Q�O:#���G�12Yb�Xns�;Y�%FW9�;�K�AZ� 2�?��b>v�m)��pu���̻L�T�O�����d�@ ����uӝo�e��NiЈ혶�CCZ���-�j;y�VN��E8Od&�,�����>@>A�d(�xdi� @�����+�D��m���և8���W�$����T8��y�#�!$�����.��:]�(�Oɪ^�J���t��c��4�)��e&S�GV4�j(j��8�p[��#`����G��	Z����%]���_q�C�%(�c��Q)+����<�2�Vd��YF0�b^3˞�n�{�ĎC�72�.���?���&ES�8'	���^�(%��Q3��T��k�$m��Y
n�,����!�Y��$����<���w�o�&��t`ײ��
�pQ��G��.^
X[�F���g��vۺ,đ�F�[_�bN��3�oݒw42|v;��'h�2�Zk�E+tu*�G�/��ܗ������/��"�f.KA3��57�3�����Vk���`�q�=�Dot��b_8�h�ڮ��� }�r�4�R$ 'Eq&<FS�w秣-�����Va�@����͵�S-�Q���ӧf�����uR��nI��[Hq����1>�bHJ�6͊������@~.�F�$�w Ei�A��M�����//X��S͢
2$/!�m)N7�h�^o�P�������Ef���TA��i±�ҵ$�
�N2�{d�e_Bհ� �TV�A'�(��iA���cU��'�������M�h��M�d� 4�8{�ׂ����d��S1��_�;,]o����<g��g��?�G�6V-��c�,�5�Q�n��A6Y�.��S+?0[u�#o��ͥ���q��@yS��T���|s��|�y��_b^�sI��;'���DfI@d	��ሼ4�Pz&菱Ԥ
�x����b�9���4�t���F��1�j^���洮�*�XO��e�#Nol�4u
��ߞRТqh|T-BDq1ir0�>_R�|���ӷ��)9;W�n4��v�r�a�npv8qۻC/}�
����!�W�aS��C���}�d�h�5 ڽZ�PR:R鸩1�Mn��P�o���v�y_���d��N#����oe���&J5%?��A������!k8��"��;��s��ρV�\�}��!X5<�R���<Rt�X�3�O$vx�b�x�e%1]
# t������[��J�(��Lrӫo��&��BV�����^~w2Λ3���҄����P@S�c�7��m�4Y�BS�gJ�P@���	�┱A/ޱ�+Ҥ�A}l2=�)^�"��D�vڟ$!�,�U�o\�]Gm�B��k�]�`#>_h6����?�J��B�g;A*����z9��\�wW���RV��u�[��Ұa&����?��GC�s����B�l�s�$�7)>�-;B��s��p!���;�`o�l@[GM���]\��y,Y矋����cr�ш��f��=U���P'��K���!�����ӡLù�]g
�O��6��$�-�&g},Z7$US]�3K3@@��b��x�_�m�
C��D�52�5�zsܹ�revR">�aً���3),�SvQt~I�KX`�n��Q�������ך�ˢx�O�P��j���=	fK���-�;T]�� ��2�RH��Tc�ɨ
_�o�k^��S�6�'U��@�AB<3r�6��U�&ow}�Y��թ !�.�����-��.�.!�1��=�ݴ~~BO�\9�Qw�Q�z�6���˕�+o^�����]*���9cgƩJ�n@ʽ���*� ��n`��@\�J^�Y��H�����$��(�
sKߨ)�b�����J��ފpU��)����f&�/R���}��ٔ�`!'����Ꮘ��rr��梷Бg�Q�� ��ॗyϽ��$�8p[��^ϸ1d;�o㽎sP�n�P��e� �h�D��8����uR����I�)Gv6���.(/�xy��u�[v���MRX�yWk��2�)E~%�Ko��5���g�le/�4�h����}��.�o4�"��h bD��S�*���"�O	��Ju�aR0}�ȑNDw�"[�V;%����I�Kq�@V����&��fԚ9�n���v��Ʌ�v�:Tj��W��	�y.v��9H��mF���Gس�S�?˗�j�����o;��R�X1�Q>c��cG�{�!Zs7Ì�=N��D
��W���f�n��0���+�T��V��N�f>X-t-���'����:w٥~#~"��6� ���eIP�u31:D_�-DL�]L��؋��Vt�����{���i���	�NFcA����)]�j��浞�V�1��*ܾ�c@%�q�)��bDCn��n����nʏ���2�����/��૒ c�:�m�Y�ޟm������]�0���F1,�Gƾ��{AqyAWN���cw%�!�dCuB�����&Z��?�X��§��Z��u���K������4i�p���`�>Ķ�lC�ަD���v}��)�:�������F�E;{l	o���������-j�iB�3�7�x8��tT&� �'F����q[�x�ʍ�U
դ�I�K垁E	 };�v8Ñ����P�s C�f	p�"4�J�U8L X�+��Y =��m�t�����U��f'��_�
W��"}�}9�����������,���}v<{�7��4j���L!��Z-�@����Jz~�/X�8��?b�y��w&C*�=2:�����;���]�>h	�@��'C��y`bUl駷���
u�jy8py�WA{�	�g�~lp�[螭Ԗ�Y?�.F}}f�>��6�բ� YY��xfs�2lxM��c�kF�ٺ~����q�9�zQ#�`��چi� }U�e���nN�xMv�9�r����k����ϕ���"ZM�{W�s�4ɿ%1V6�.� [�}�f]����DG1K"�+6�܊�S#e !5k�&,����>��-�V$x�A+��к�8���ci|����ڃ�-e+������,��X�^�O���2����OǟfFD�MZ@�3=�'K���2M�s�z��Ԃ���M/����&
A��:�"!�j�B9��B�K�mѝ�7�N�l��y1Mdh~���ֲe wj�w&��"�^p�4��\�F������6PņR(}�7Ba����,�@)Ω����`�o������_C��5[#��=f�<�Z0�	KA����Y�Q�)�+ =��	�ʐ��Uݭ�f�2��z�Iى�3�I�mNs{����lɸ��p�p=$X�l�Zq����Ch*�L8^�Ff��W �ȩ�\g�����j���?�T��?�ֵvb ��1�pHO�I�HJ�Z�]@��rO2�:��%��En�����������(�o��p���6�F�&pN�����J�|ˍ��%�Ϋz�+�m2��zaO�Wa��A�/���ҧ&�|��-�/x�з&��r]z�>$%}�?�?�n��s�*2߽���{��0����9/j�_G0��|p�=�6���Q/6hUe��	J������8?����C�Tҍ��"!0oFR�(���T) Aq��{����k�;���05����w"蕍g���f�������PX��<�c_(�\?N"��qEJ����s�>ȗ4���mk��x���(�r�%��Y�Ki䋑H����)�_��;<��+��Miy
�c�s�׏�󷺚ڪ}fk�&PQ�vǤ��3K�_�Rf=ʟz��/��i�̧�T��{���WdSZ����<3\)�4�?��[t��pSL+_0J���l�f���3��#"��w�%�B�[Piv�& �����E��j!넻�$��Qz0�o/��F3K��=����6gdoҴ�۵��20�{7���!��PU�p��։����*��x�:��
SD�a6!�r�@�W5O΄�@��wA]��0��b�}&V�lL�|$z�;y@p�)N6V8�w�cjxw��]G���<R����)�Q��9QÞ4��7��E��)>�KM���@����z,n���c��#�'|�+�W��.�ٔ��Pv4s����t�dEYB��L�]zi�k/�wa�i�OO���bL�i�+��T���6�o=���q�^�p�h&2��1/Oװ��\Q��q��V|��|)|�G���q�pw5�7ބ{^�p8C�sсvM�K$vqG/.���p��0�(��AC��L��d��^�9	wQH�1�u����/�"5̴��1���D�w׀��Q�]�@k�dC��J��=fǥX��:{}1Fs�	���o���,���L���p�D�|+�b*h�p;�Tn�
6jZ��'y6G#�y�vqS�*�{��,߷�D7�Y92:�Cg"f�Z���>�����'2����?-�=���i��^Htۚ.t]dT^y��>����ڽ�H�$�����a���K���$#j�V����/�]Z�yX'���; ��1f3'.#MP_f�Y�f�z�+ �C[�!��~7����T���R�C�4��f��Q��WB*����╇ �9�mR�xI�b::d��+(x{�_��0]Oy�U{��,�VT���5#�o��+�~L$��<�PE��M5�m�#��q�[^�͔�(���icYj�1�oe�v���*�wG�'��KE�m8�
�吇��� S5���	���?�ٻv�!�{�i�)��ncqK{1e𙾨��W�\?~H]�j>B�M$���������-=�̧���]ھ�W������X`���m�
�O��mҡ�+j9$c�j�Cp���	4ѓ&��4�2'���R�5Ⱆ��2sl��h�n�`A�9��P�JW�Q�R������g�/-a��.��r�ta��o�C}�f��{$7ϟ�?��q�ך��'�E샒#�'$d������T�m���=ܴ�&�� /�9^��.2hV=8ln��O��$�'ř��M"�>���( ڬ2h�u=���O�<�wZR��1���L���!�i�\���
*q/Y��p��68(��P�)������R���x�_��������aYtߪ���%�{���=pݪ��7`�01?]0"+�~�_�a�\901��,���DИ�������1rUQ��t~�3ZQ4�_��!g�
Ħ��b�9C�5S�ќ���� ����N]E��\���V�$Q��'�" �e� 5�[�NT�G\4NG�{�����~�dB@V��zŴv�ƅ���*B�vSzM/]�oq�8�m\�JW�T0.����m%��h���p]��l�%�)�1$=�[�)XP������Ƞ����T@���，{�5|	�y쮃+eJ��?�eP��v��c�I,�Ma�yN�LU�;���ߐfy�2��h��m6�ۃX5\k9R�%��8U�_���{�t����8��U1�l{��^ ы�Cd7��m�6u�����Dv�g0b��'&L�Z:d.5�)�,,�d;�2�Fw\]��Y ��`�����f��e�q��ޡ��������Z���EN�O(&�C|������w�v�R�����6PՈ�&&������L��ڛ�"���A\nxp�99�����I�:��}�:�cP@��;pD%�#Mu�;<��N
��،�pT�����.1^�O��$��0��$�j��4��RS'�U.�&` a1��a_�հom43 raPd��=�
q"�QͿ{Wч��P|���-�p�����@������v3�y6x��D4ye�R��ke��I{�����L���u,6g��W�:�a8M�<Jzq.���i��T��x!�	$w���QH�/Ò���ˀBB���������ɏ۬U�u�{k�)��VZ���n���j��"��Sw`�5��,������Q�1�T����2�SH6ỞP�fpө&/H��Y�F.����52m�$�6ЏO��<]��t�E��k'Gsi����������`Ƿ�/.�0U�&����B�?����8L>�DNI�}-q����d�ʀ���}(�g ϶�K�N��i%C�`��=��s�Q��RXh��W
Ά�aR���%��_�@�扳8������}��V�c�x��BH��?��c��Q�ɹ��b���AL�:_��f�Y4�$�q�{�QҞ1��7�	����L���ag�j���Y�N	M�.C2��>JO��(*�Ϳ�:�ԝW0P�����{���+Z�t�)zM.���`5�B=���d��?m8��g�Q�!ێ��Q�e��!�z?��ӽA�����<@P��A�^"�e���/G�d�i�����aI*C���g��s�<jo���}��h`�
nh1.M8/�Rl�
����y���Y!�C=p������W��T̰À�������R̰���
��ia���+�$g�͐C,���q��Q�����I����.A������s�B�0\�d�#�7��#���TI�Q���4[�37�7$p��	.�/xu�|�v����r���M_!l*_E�����X�h��%!HB���d�?`
g�'�ea㻄ʰl�q_�kcbHX3�b��m��B���4?r(���:w�oe���HB���|jyAĲ�gi�d�as]w�?�[���5�e� 
[do^r��R���{�/�����.�&�ɓ�[��΢�dY�]A����Ed�/<+�b�#��(��뎫g�V�'W�rt �26q�jVҟ���A�`��V����T���`�̻7��ә]&ׯ�#���^�է�{G��oK¸C����ۼ(�
�-��G`����8Fܨ�[3+�3��(�i���D?밿�j�_��
���vz���f�㨕�È�o�o ��B� o(��y��z	/���������MԔv/�Pn�9��: |949�Ӭ���Y[}<�<�V���0��r�b����v�H�!GQ ����q�ע�2.T��X���6u-h9����l��'��GL�8�2���'�r�H4N<E
?����|��πJ�$�)��=�/WɟD�@����]3�\���^��T�j�m7��;_��1���؝F�.�D�Nc��G%����v��9����1���x#�l)��-���^򳏤����}����MU��Wh�U��y���D�7���#I�{k�uz�7amz�nl@Մkkk~������C�a���C�DQD=Ŝ^�'e����j�7[�Э�c��[}�e=�͉���F�K���%�Lv�{pQ.��X��e�HQ:�3��������b�+Mȵ�[}���v���VV�#5�8gֵg!�W�m��U6Z�B��]�С�v��ꆴ���c��h��	�@쿅% �u-{�P��@+ɔ�F�<]�T�B\H"���0�e�H|;��YYo2'+�<c��\�t�Fm��l��հϬ�s�)]\R_�Gy7�2v4��'S�������6��z<P��ث{/��,�n�G���/�L����K��ʢ��X��a�����:,vG5�_��9�R�|��ӹn}��������h��>��
D�E�4O$N�dj��R9Jo=p+��.P�������{BKϤ�ꐛ�kC��6�d*��kQ�H<$.�l*5o��|���(��BT�4�+\��$Y�E�*O�i��I*�u��?t��^l���3��#ا[z�1J��$HO���0A�K���\G]T�I����K��Y�ٻ����`<�|�؃b~�3�7����@]��=�6JͺɃ��ĮhL����������'@�x�%Ud\��%P���E��#j��	�n����ё,nB`$[,6/����[�!� �N�r�0&oڵ�T�
�<p%ը!y�kl
VV|�o`D���vm�}�ʈ���Ʃ��̳��u��,��V�F:^ѯ��G����]mt��3��r�>B�X���!*��%o�E=�7y�@�F^�֤}'#��W���lH�	��p�3!�|�IX$��x�L�VZ����d�:���`��.�ጅ?W �y7�2����cg�����ClG����A�:��4�|8��~bBZ�\��C�#�5�m'!E��7����������|�l�d�ڱ�Ro5-�����#hǟ��M�Fys��I���4�������MC^�^ͼx�\׎���pS�����ą��3i#��h��=�9��?
yX�Wmb�ɓ��|��#�vrd�����8Id�z��Fh,�b�-ܲ]-ĕ[�:��_.4�AZ.g�K�m9$��3�!�ߡ�]�2��s������{5½I�X�W����UT`sLQ�}���H�\���:�[V�=�c|(�kR�fu��ޭ��}�M$1i	,*�P�(T̘?gQ՗�"�m�}:S�A���¿-3���ŉW���6P�8��W�4��a�oD%w�S>���l6f���q�r�[�}����n�i|�VG��@���-?��ɔ��<�p��"J���a\ϳ����IB}�0��/�kr�L#A�m�'�!�'���BX^ˆ����6�Y���q�ei��P���a�\Ğ�d���h縭p�G�KO(z�����]��_��[M�XT�gͭ�_���W�C>oT+�U3��>UE�!��x+��3�qf�啦Ð��X�Xs큔-����;��&�k�|�^7c=�dP^����t)��§�;V����4�:}��8h��x�I���lw]�T տg}�'����4��KV�o�F�u��޴o�0�,F��_'Z^�� r ?g#nE���y��cJ�)��9sI6o���G�.U�Ϲ&A�1���s�ʃ��rq�J�Vl	YH�棎��L��R�#h�?Hr�I>�PN��p��`����&��o�6�ce� ��p���Po)�Xwt���yl5W��Z��צ��6��J�T 'ql:��m+;��8|U�ȰЉ�h��=�k$9�?`��tW Uq!`Y[K�~�?�7$�9�_Hb�w��H?�|;�΍!�9;\���?R��
�������O��Rz
Ʌ��{��=���-H@O��y.6<���(Ų��$P1ͭ��7	K�w��i�*��I�g�4�k�?3�8��ɹ:��a�����:���
0���9��7�m8if�[U�$M
>V���,�Jᆞ(�ȁ�֨�� h�W7��N���ߢ�v�S�5�$ё�J�gƍ�44YNI��VdÉ?A5��wN�,:_	��/OA@����%@C/�/]�a�N�*�ݏ�&jA�8,�@	�a@��I�Ud���SMT;�F�5��U!Q]k��S�#@Ub�,����i�g?C����r	K��_t�>1,{D }T�楮ܬP��T�{�Ѽ��gW~�߅�o��L�� ���Q�I��#d����8j��:�)O�g�F�a�'�~WX@RV�Bp�1���Sg�|I@5`���Tg�z��	�Y��B)��|v`eU�����kC�r����pz�e|/C,�p�x�c���`r����P����)~��o�>;�����#�$�d�ﳼb��rX����M�ɫ3������3A�Egl!� 9k&~P�^H5�J��A���PsF�j����)��3hJ랢zb̕HK�L��}9��d��6�wr �g`���t_��؎�b$���S|�ā���6��W���@D�օ˫5��F��x�S���H
y0M�dm����Eԏ8#3|�-���������Kk���%�~<(�X��'��W�Ȯ�-ߞ�p7cb���c^W���0(�r���o����V"cI��_�_�)���FƼ������ޖ�U\�&���1K����Y�����zb����uF��j��x����Qit5�����(7U�n$^� >J�6�R�������5�5���^��ƃ����L�mڭٸ.�� #�PEX��Μ1Ƴ�z��SB����-M���ԭ�G;%t�*2o)�?�("�tf�g�0�h
�:r�+����^�H{���2!Y�A�7�����G�J= D��;o��K[@��e��5B}58_�i�Ń��E�`�{5�ZZ<���H:I����/�S�Ks%�T2����ka�u̤c�@�:�7��N2^�'�����P۟���1���\����q
��4וԊ�[(8�m�Nn�KT&fu���G�̈&�b�	�R(Gi'mTѺQ�v�
�_��(�nֈ�"��I����u�/�.+�?��q�kKmYf�bi�8�S����aWE��?��1㫧�*���w�~�\ⷍ�"���P�H�8��D�Tu��,�$�#���[�Z��Iq�������H�� Ÿikz�1�<�_i�[�c����e�#�l|�X�Qg�=# j3bQu��ߍ�(��k굥�5ݔ�~~X�e�j�u��rV�pl��)�8@�.�J1�!�~�v����y;;��<^�#�k�3yj��
�6Ȑ��2�����:�Q@[DA�T�D��i��Ⱥz��%��iT��N�;�M%���Ҵ��W�r�φ)Ә4ĺ��rS@����U�[C߱_��R��U��ڪ�|Q�?��3*7��]�;L+c�+��h�/t+�|U�����a)p�%��r��n���;���Kt�R�Lb�hh5Af��#�e8h�f�)$ӱMK4�Mb�)zU�� ���_F]������V�^��ZqV]2^��/+����W:!)E�*_���I9��'��KXZ��i��4�o���p���OO[��;��kH�u����[�>��`<����z�7}���}qG��z,t�8�B俑�������Ǒ �%]�7>��I�^��{̥�M|5��B��6ʱs��cH��썯��>��ǣ����~��s�M����1I�V�]$�>t���X�y��Q�<&&�$�j�R9�~�w����������q�	�V +��)A���}������ �j�D�(�s�?n���RKPy���5g�HHY-tdv#�^6ڦ��S_�yx��N���k�I��	�wg@ا"�U;�/���g�e]v4U*�V�v��$���q��<4D��:�U�k4�F��¹�(m�t�/���)��O��?7}���JU�>sk�:�ൊ�jn;�K��?ꋲNZ���!���q���4~���U-
�\U�e�a �Ibv�����g����	P� `�b�K���Nn���8��:].�,�!S�����ѝȭ��ɥ�E)�f<e�8}�Tƙ��cP�E������~�	���K��%��:��*�ܓdC���X������ÿ02(�]�e�����4���W����rA�ܐ����-�+fzb5(�l79 ?�9��@)�� �qtT��R	Ϗi���=�~T�!C��
O�ΝS�Ż	Dr�WWpw�����wm�|�Gem��&$a���ҥyq�>6���xy���]����g��;�EY�O~�co@����
�E9g?G�Q � H�ٖͨԑQ2��]T3{Q~��;n0?/��^�{��	�{�õ�3Gw$V��w�
�24MU}
�`A�)��]y:��XφI�
l��M��x�wI��u���� �Pˆ�q�>�s�i���A�#�3�ѩ�c�uԽ}K�zJ�E>�'�5�]^-��5�S&��� ̧���ƶd�Idٻ��Kd~G(~B�p�8�q���J��'ߖiYTL˝辌�E8�r?:? 6��kK��d���N���1̬���,��3�!=��~�>CV��H����a�������:��YR?��68��_�ʥU�5�Ϊ�G����a���!)�2@M�4���;�����Y����&u��?�����/H�,5���\dm��s���.�K�q�[��y79֮��7C�6�H�lէ�[��rzQa9��Ƹ�N������C��ӟGǨ�u��̘a�/��*e^(V�mF<�jƁ��G/=T$�dagk]�h#�b�j��q� {���<V�h7}��'~z�LM��"4�1`ѹ��
��Q�ao���Ff��߂_��.kd���z��!�R@;�|8ɤ�M��L���+c\cs���r.�⩦e��7��&L*�4a��O60���~�,?����.2/]o�5X�s6'���F�����6���ڬ�wO����*GI�"�p���"Gf	�=�� ��L��1V�����;W#1?g�^���s��i�n����T`�`m��!^j�
�νSV3oG����E<>�ta`�����}�2�Aֹ�SŽJf���D�G,|��ˤV�eϯT�	$\�S���ʁsnQ{)��ۀ�d�23��mꛅ^.eR���ob�ؔU�6�m#!�ZScՇRκQߪ���E�|���4��T�fm�v��=�CN3��N8��7X����~w��I�w)bk��R[�����ʢ.Z�.U��h��ka�\��U"�:�N�ZD��;6σ|�_ȉz�	�ikvN{�TYL�>������<Q=M��Va�\(�N�#�9�|]N�K%۴{��U4�&�Y����'���7�Z�u9u�����o�x>���9ͼ6��H w�Z���B&�tڒ�^�A����ه�>�pAD��ݏx�K��\�s�y��d<|5~F�$.QSS%�E�_A���# 2���|��!�bɄ���n�,��;��3|�M�q�`l�X͏+V��A�+*�C<�'C�`'I������)襔A���]�9��FR�j虯Q{�ed��ݺ�:�#�\���uc�6�e����(}6��Yʬ��h@�߭�T_�J9�)�3�F���R���4���/�>D�`��h�٧�	�Z$U͋��U�n�?�߉��D�Z�)�lH�)лg!/en	c���$�f|���M�i7�4��� h�8���#QFm W�mz���/�}���H�S�
��y~�qL�{�Iǳ�S4O N�y�Ĥ��6�P��B��.Gy��C,�]�*���7>\$��3q�G�cvu��C��:�A���R�i�:v��@�Kt9Ñ{�����H���M�����{���%��_>Rg�멼@���չkN���➨���z�g՛�i/���`ܹ�+.B,h�:�l� �٦��ܮ�+��㤪��UYwIl	�kݽ�����ue�T�r����w
<�� �|����p�o���;�]b���B	3\)�ɤ��V$�t9�/":�Y/��+��G3g���*-��}�P@uBU\�U@V%��͠!D�lk�50��@��ó!���'�5l�>�u��ՓxX�4v��zp���zZ��ȋ�r�뗫d��9΄��l-����(�����o��7��
~�m� 㿡�oU���
�� ��~iB������%_�u�����7�WA��S�в�T��)��w�cb�/�d�M��R+I��i�q��55�27ѓ�h��L�!qv��t`����Ŋ���O�~�3*}�úN����H��'�8������p>�2)T�nK��� �U.;��i�-M6��Ga���N^o\1!�㯆��m���~�2 �+� ���M6!(ݓ9\�MlS+����()?�$_vJzyvы�����I�Bf=��#�SIM�� d�B=��iv.�)4���˺��� ��@E��Wn|i�w��V�!��]�Η��Z=������F�z���<?���!d��T�FP�ffV���.Z)^$���e��	�x�>�t��H��!a4}�%D�/�����9v|����>�
0bw`)��j�p�(H��dbN��5��ڕ�(�h"��~���:�G�$;ܔWN���?���3 ��S>rP��>���}����퉆=��#�' f�L��]4�Lhx܉���u��BA}�͜Q��n���B��FM��9������Q}G��Y���7���g�#bv���C�?E>\�� w��+�K�%2��ͨ+�y�����Ƈ��J�)���{=BS������JTWT�`��5�0R^���1�1:���|��g�ů�����>�����b�T)��ĞlRF�[szK����H��H��$U��n淅Z��;�����9E�lQxZ�~���1�j<��Ҫ�
�4U��3�X��?��ޙ��1��g:��f�UCZ�\�qu"In�SWT�-�V���K�-M5��Y�8����/uh������[�����Y�a�?V����B�2JnՈ\w�/9D�t������S�wcp�E-/�mN�A�����T>�'���'�X)�Y���i˔�4w�=1_T��P�PM�����Ψ��=gܩ��l��د�X��2�(Gত��H��0^��E�8�X�K�N r'�YǉG 6�D�{@��:W����6.#�͟3�+���eT�4���TJ4�G�*>��/s�gOɹe�k8�g�E�v`��ae�R�_u�Ѫ0usk�0����0
I�F<.�^?�.>��A�o�1ermV�^�XU��� ��.i�\\��Іl"�����^^�yR���S�c��f����*D	�9ںS%��s�2��e.��$�*)��#�Q�Xq���a�c�l������U!�����L�f��?܅��~�IOP�'���u���>�KQ��mh�c�{U�ѽ�Ip�]9嫞�8m�'DB�!�:��s�5��}�W�up�q�y�D����}��B�	�-�t�7��	�}�b]V�F^�c�}�<.m���<���������C�qC�b� >EhŶV��N��b�B��19C�1��F���X��6�Te\���(ܐ���s@�nKcg�o`pi�u�lm ����D�ҔBE�.u��L�!���!{8����^�zB�L��ͫ�iLf$�Y0�H�c���L��@rFNp�@�B���E��I��*T���4`U����DAs�V2,E��"��=|�I�)�JcJ.�*�v#���U�w�3J ���\��Ɛ��������m�m��!DF��
;"g�wvgnLv�g��=d�c�S��(�q����䑽���q9b�K�&Y�k=8AQ�|$9�쫥P����uq�� z|�-��OA[M�����5î����Ac��+6��JI�����r�=��Fsn�PP�ŨA���F��A�n�2��r���e�d�xU�Ak�i���l���e0�^�[�����3L=��� "�j2O����7)�J��w�>�:^���C�l)�[�mk�������m���(��s��,��_e�6��E�6UeCg��M����a��µ�d�������Q<u��La�a�'k�(%�'�P��,�T��]>�����Ƴ��7a�"��Kv��:�Ǽ��h$��n���R+���a/�:  Nڈ�e vF�L?�����c�`�`�N�!��)>8�u�O��0^b�["�x��S�G-�ڽ���w4�� �oe�b����邈�'f��<2����� o3
d@��z����2�ee�U#�}�§��]���/$&f�w4�S�sI��0.�Q�
x�C�<o���;PʑRd~���͠s�#� �{�X�3Ee7�C��f�7}�Z��a���m��`M�B�ֶ�rfZ����r��b�3N��)	�n��d��V��zq���>E�]�����l�$�L� �^��}�ơ�R��j�{T&�?]��hk�"����M����0-���j�{,��[~AW����f���;[�5fJ�\�"�%�FD�:yө,T��H,8��Wm[i�mk���l�rw��Qg��������cqn��SN�dГgM.�� I��^Ju�!j�;��R>m,�PB��%�4��5�p-@�ɟ1i��@f�V;t&F�����A���l��1[�/'���">i�W.�_ p�y�� k�D���%O�C����j�c�t��؄	7� ���7�O�9���Ds�[���T};�,����,�����9���%� ��K�/�r@͠ Yħk�2�>&�t
�j5 �Y)|�x�Tr��=�(&��5�hBFy;k�-�̠�<��E �C���b�P����H���<B�*&X�H�<Ruأ@ �bќT\3Fc9{PBM1,���[��\�I��t�͗��Z����� �J˿��B��}ȦH&�F�3��*Sl1{�'�"�S;S\�~��<� |J�A�W;�:^�8<�a6
�7O?�g��jo\Q=�e�ä&����>�n���q�g��&g��\�Zx��:#\[�����1�s/�NV�Y�.$��{��4��#6˷�j�"��niw�-��GKh����VʂE��i#�;�����kI�fu��A�T=�4A߆7�Tf�pN��a98&HIε����ʫ�)A
c��<�HO^ nRޗ0�,�=n��͘��y��4��#|����g)����զt�O���yv
@`
�C�"���c��7�5��+N@�/t?� +���gc��ڙ�1I�D���ˎ�l'����z��H9�]�?�GR!���� ׎�2t�{Y1�g4*�VpVd�{IW���HȡXM�E�?i{�<d���ǋz�S�yQ�(��:����Tى�9)GLBq��]/�ϖE���fԆ���ax�[�wK��P��*���a���8jm2������������#jw������u��c�z	��"���P���Iʺ���1D�̮l��,�r�et&b��7����:Z��V+���׷{>�>Z��Z�����F�;T�`��(z�,Vկ���^/㸺��#���'r4T���$B�n��Bݭa�`�=����#D۲�9�J5�2�G/��.FԦ�-���Z���0�P���g�#�^�2s��C���	�Z��P�R����]P悑�4m2d��?MwZp;	���8I��~x������[���{lY�i��;E�G���T9(��I�s��
?��PRJz
m���<���6/���m��`����nQ��h�8i�>B��.��nC-~�������~�貕����"VG-?n�w$x�}�Xen]�3Q=K�Vx�%��P��J�8Y���ʏ�OZr�Ow�_�*��t� �8�b많�ˑ��~�
�yb��ԙxo�n�-�� �z�u���K������:��|n>T¥�\�ht	���kx���
�Y�@zVt!��p��%�u�����H�؅��z���[ﱡl�a`I��'��6�q������ȒCh�I��f�,@%����b6ע����뀰͡�����/�TO�y#4ӟx�9�LP�g�(k�Ν�5�����z�^��Yry�Ik���)�:���H_yIip�hIHE�ʛ^� �p�)?�8��Mt�����a���[��*�>
ӟ$&�r$k�N���_������x���x���- �3��\\2��ׅ�H��W�K�{�gtL:"�^z�>{�e�7%U�@�F�������������b����0��zB �a�XW��I[�v�l�?�m����;�J�{�#Id����HY�u�9�_8����,�B_�)��
�2�����-)̯��h[��F�\m�WΈ�Ѱ��o���^����c���\��@�Of�i�o�k��ݗ��X:�e>B!U�LM'��a�&K�CCd�U����9؈$Pi\��
�/�~K����_��Q������|�eɓ�t�eD��h��
����}���)Zj߰�w���3l+׼,<����0�m��<���oN�59u���!��-�>,D�tm�"�N�7��⽋]�-���H$�&x�]�qD6CAWr1��^��L����3�Ȭ-ڴb���ԡ?C����~ǡ�*C��L��)�?i�g��M�e��KG\r7�d���i5�?�\�N�L�x�s�W�9�q��"��s��?J��d�7Uu�G�{r?�����ܲ�s��T�M�k5�93v��$��W�����-G�m  TB�n����+��@���<�' �:]N`�����6f��H}���l�*A�u�Y�W�E�4z�"1����y����\;D�Y�|�O<�� ����(��5%�Z�R�̴%��3�w��>��bC����߱���+7=�Jl���l8,��|�Pa�Ʌn�:`) ��l��"���B�_ؚ]�U�G8Ò7�?(	�@�ބ��a�a���{�s0�ω�-+F��y��_s�8I�D�Y��U�f�>������"��x���B!��tjQ��\��A�p� �y#�H.���|(�h݄,Jȸַ>&z�.nƛ�7�5.��;�2����{����c��˨�ŴPo��*�.����e~�G6�v�o�\�xb�,: ��%0�K~ ;"L�:B*o�k�wvcʯ�І�L�� 1�e�
c]]�����C
f&t̺\�%�lF�qq�"����k/�<U�A��z(�7���^�`�#ro�dy@)w�mM�K}3!�4��䖥{�_g�D�rǌ�����V: &�Pk5o����Lw��چHq��Q��� �N�i�J�2�o�vS�K�g��5�v;{P07VA�p^޾!h���6AA��I�(l�	����HZ���J��2�+`[�L�-�)���Ś���wo����@bA��h��cv�Jk�V������s�i͆�&|�nE��䥙��
,�����
�Z�]2��R�tY,���t��;i��{4��s\53�pE�"eZS��vH#&�]�,fgȄ&a�iVS|�2��ZmA��-2�:�[���	x56͏����2	��D&�o;$$��w���E����4$ۥ����/�����%�OE-S�]�#^lg�zd������>�yt���6l{f�-�#i��-E�#vJy�k�˟�œk%�j��!����-Q�����HQ�<����eV���Kq�K	�]�I��$�e�$'�q:�-�UhBz��D�vZ�D������%�2�fѦ��ɥ���EPpƣ�	��p�W��>Ʋ����Tx��̊Ttw��LI�!��B�`@Kh��[YkY����3��_n�.�l&_iCd�Iw\<�B��� �Ƴ���6�&H�죗h�;ː����c���5�Tu�} [k-�Dh�� �QAA�J�yVtMU%GR���cM��� �Z�X� 8뺭��o��%s���r�*��}:�)"�C	���U���}q4�c�_�(������64���	�w�zy����>����,F�ߋS�5� |X,'�\��P����ExZ��K��2^��b�O�������ݰ�ԧ�]�	��^5�����o{�.z7��Q�J�����|�w��h�޶��L"����d�F٦��e�/�@�%��;�l�3]�l���w��YfK�'c~����9~mmM��Q�3]�Nu��=�%�3uZ��.��<�x�0x������y���뚯���a֩�1��Y7�E��T���W�6-����M��0�
��ucOu�ʨl��6�F��|�rD���@�l�G��.G�I�v�!=e(Y��oT��	c�����Ċ��EÈ�����(	6d�k�rފ�CC�L�|">~�����+`��%�O�=a�O�ljm���ʓ�'�Ƅ��|�b/Ƚz��q��3�M¶P [�.���X,��m7�����Ɗ>�NAap	+�3CP����_D;b�A4հ�"۔�lW��_"����^�`a���^F]�������J `c���J(�_����UF��JI�C�\���� 3H��tO�c\Tbι�Q?*%J?�&���D�i��������z&�$��AI1 �r�� F_��@:y����+��`9�R�b��FښD���|e��e�χ� 3����٠q�N� ��hkT_]3����Wˡf�ZG���Z��.4fe&���Ȗy'��M�e��Ո��?X�Fm8rl6�|��2�v�?�?�:��Q����ga��!�<бp���l�<o]��$���M���jc��a�3���<Ck����-q��P/>���|��<�@+�x�P�07*�RŠhV#D{V�x�7󽮔�xiE���S�����=�n�L	/�f (C{�@\�H³��@"�ߗF#��I��;�އ�O�P�p;�F��,�m
C�K���_��ЩNkv��� 9h_C���7s$�څ�}5q٦�@��l9�"��W�HAz�j{�J~2��:��r�q4 ��؝�:q��&�:@�T����;�}�5_��K��z�����r��="�����Z�C���l����gI�=����1#�����9n����i{#<�	����d�?j��&,�`����y|1Ԝ4�kn�f����m�S�%�CmG��2M��8����~�g�3�L$�dF�ho�z�+�r7���<ɼ��p�
��'�k��%p.�{&�➭�������IpV¸&��������K�h~�]�R\����I�e�S)���M��S���88�>�؀E�AKԖE�|�.���<T�0��2@����ďz@����ELjx���?���gbO oJ�E�9����\�B��~h�f����$T��I���W.`�F5d���U(�w�,��_򲠡1�jU�b�dGv"?�%0@}%�h��6ZNĊ��<[k"$�����[{����Z�
bΜC!�Иr)�%zJ=$YH����#�0\	�K��a�j�g۸]yp�k���{ K�@��(���0����e���K�C��fHj����ጌ� ���A>aȑ�ɜ�x!E�BlbgXʏ���rf(��4�J�C5M���SB�֥gf��� ${^<�`pQ��[оL���Uu��F�2\;��&,�J��p�zw��6��{���1�� ;�{{�m7��r���|�)<`+����t��p�FW�6�qQ�������5#�R:Iyr�eH=1�Qx-�����ְ��2�+�����m����;`�F�|�����a`�L�f�X��j�Z/��f���F���7��O��I���DЊ�Oz�v��&D}]�$�u����b-{�tȆ�� ��E���ڬ�ܲ����A��`C���	#�np@�ݭ�@�<�6x�E#����*��_N'�]l�	ȩ�n��9Ζj~n�fČC��کA\��ͻ�P5�����1-<���3%�}�O@�J��0�YA���E�d�f�%>f�w��;� rT�j	�@�s�J��W��k��)���u���.l��q?�/N�^)�Uf@{�j�����J�-&�8ɘ��Wf�����4�b�'P��?v@*�Ը��i�}��-��h�c�L��'�<\�W�����n"H�{��6�ؗ����4���N�֯�wVW��1�����k��̳#(X��1X�ar��u��:��Ӻ��) �}w��;�K�e����D�d(:0���#��]�t�񾈋PMn��N�b�m�`VeT��$��%f%���8�&Y���s�J��<���ԨpagV�s{�M�[���$��4�Ȟ+�P�I�Z���ء��ސQ!���t�mLM�'5��/ߺ�{i⺞Kȕahv!5����jK��T�o�����<3:�&�&��{�d��W�h�J���߇��]r gwr]�[q�y��FKZ����$,�y���"\��T�n��#%~�{�&���Er-!~�Y�g�
��VX=�LS5ᱝ���k*Q��'��P�1���d��q�N��F�{D�{�2A���oU������:�K�&"nO�3�<q��X�)���Λ,��:Y���ګ@?�Q6�Pj!�~8k�=ة]sv(�o?�"h$��RU%�&���tW�GGz�o1~�y���b��?��I��R���^�Q:��Vw�9r�R�pfsn	t���z�U�N�|$�0FI1ۭ3H���S��T���s�m���0��U�K��l�d���O�,�\M���մ�����>���S��ۍ�y��f��k����yH�ثe�/��δ����iSF&,����	�u�T[e9��vdBD��#`��%��Z��e�cв�;G�0���U�Ub&�t>5Rr��%uE����FqV��\3Fk�N>{[l��A�|t���*N��kJ[��}�o�c���\���ѣdX��.֕�� xh
C�կZ�%��0�$�=&�w(�V�I�Ԙ�����dX/%�1 �-oȐ�#���$�ѱ����5Tsg��B#�D��疶�� ���Ԕ���\��#�{��\ӆDZj_��3
x�<)�d=�e���+w�az��+���FV�)��U3������R^2mE���l����Si�|���%���ԭ��gү�0�G%ߍ�G�<��],�n<E@�R���-��z�p�IA�?O7���,@�]-�-���
�����91cAV�֓�5̍P79m�3�^���'��,a�x�]��0�h�9���NԆ� ��r,z;j�:vA1�8�}�Pm|��#���1e�¨�́��s;���e��z<�\�G�~E��R)b(�=��~����FU=�l�F͐LVXl&w��4����$߳/�k�i���&��MW
�Qe�ѻ:/X�=}�2��m���/��!ze��v]�R�Eh9� .x5�tӿ�b�|fC���ApcjR?H�b��E��EY������e��%*�j/�@�����P�S�g�tU6�tZ.�KU���7;�G�4���@�Uʉ�uLs:��
���WlK~�an�����e�R�9o�E����#�*�����_��gՉK��
������U]W�>�4|�T�&��� ��L	s�7ǯVD+��&���J'�)�cD�2j��(W~�&(�xA��ݍ4��+��Yj��� ��6�����[;�J 8U�kљ���X��F��0������1���'��06�U��6n:�K��r�/=M�t��zP����@Gdlv��Kr8���N�<21tYm��?�n>3�������S<�r���א�y��!-I��]�RE��ޙ{%#�b!a���1��둒��'�(��f�{�Y�W4�H��QE�� �Q�6�
ԯ�Ϻ �Di�$Y]R�n ��i�#��m�U��.��Z�&B]h���z�K���#��sv�s�Y�]�n�o���:��F94	�H/@������aD�-�߅l70��Џ�1�7��2q���i��~+id�uS�v�٨c��~��ٵVyb�{�&p����lԿ��E��9�*�)�V��yf��f+
��a���5�ϯ̉٭��{���Z�c����@{D��e6�9�Pw��i��(���}0N�5�����~�@�oW���3w�4U���D�jNի��;���㿍���{��Z�m����6|�{^��|��@�ǫ��l5o&�(�ڴ�Ԋ͙S� ?'�#�/�F�Ag?@�����O�o��Z1�A��^��wq���Ce�v.AdsQn�PA{���r矪�S2��\�O�b���ꀉz]�'�1��@����IA#$e�h��Lkek�)�����RW�����D >?e��uq���ٿ�m��%d׍���Eݑݢ�!����\���M?���o�)�ǿ$.ō^غne1�w0�xH�~�z@�6g�b
t\�ج{Ȳ���a2Wf��04�E`�� z �ʐ-�t4�5��I�p
�L�g���u��h�IX;s_{��ƽ���o_S|.��L�]�\���;�Z��נּ��d,F��:���gL�]��23$�C��b��b2��wf-	~���(K��*�ʏ�=@�g'�s_�&�ȇȴc�]�Y=	��.jUr����J���Oա,~�hh���H��6���N��e�YB�A�#�E3U���3�7�'�'슟ߝP*��Y�K,�M�/O���Y���g d��Wd>�b����4D1H2�C�m�rɘ����f�Z�,��d`D��禢N�g�n)�`C�	�+��{h��#*'�e��ډiP��iiLp�-���������	:�j��nc��,Z��t+����R�}���t�\��������TZ��FДD��H���^�����8�����$�צ�]�NE-��j�_G�D�M(8
ڬH�Q쎀4�yx�𹋏�Ě,�1H���R ��"k(
�b`L���s2�������l��X<�.��xƅ�;X��ir_��:A��*�|�Q�#�j�I�{~�TZ�� �B�nA�ŗ�,�狞(�����}�k =�TT>�|q����cYO�r ��?�� _�{�)�������D�p;��8Mul���~$�҆{F���'�����oP_�U|(��P���6�ڊ^��ֈ�(���|���M�kO�G�T�(�R�ϩ�ڞfl�*���O�����3����4��P�jQ>�����HK�e�_�3�[]^��i;�F1��y��'��ef��F�BW�ίks�X؁_M0S�A��ѹ�*���=A!#C�%�k��{q�R_T�k�Kc��+��>�wB[��iM�� lZ*�o��x�;?)���џ�0zy��!ޓB����_�5'��`ϾA/�������c["���M��mR������e��snN�$���	��O��LE\�^
�8��
��p�0V5�_�e��:A�0-�t�|�Ƽ�c��Dh)�8XO�RrB3c�^���-�7d��N�jP��%ĳ�B%��ut�6���!����z���G�U�|4�Tëڄ�e�V��F�m�"���}���\�5�D}���1��z���������~u���@h���.1-ۭ�����,�Ӣ?�!�%�u��xnT�5�?��7kb^R��jD�-�t� �"�2aб��9���O�Xܨ�1�V�*�=fO��֜G�O���\}Ƙ�(`E|�����x
�cp�X�#�`���!Ұ��T�8,D���~<UH��+I���f�"�xM���R𸘿f�����.�Й>T�>u���x3 ��� ȥS��8m�_Iw:6n3?�:�����|*#�<���tM��& 5/�����ߵ
��ڸ�̵2��PJ�����>IO���	������
%�ˡ�����3̋N�WXB5ղW�H�<���ַ��4	#�)	��n��P|��٪�"�vru<��ﶚ�$U����2�T2�s���'��ɢ�E+th�.�TM��C��ӭ��_�֪���q����f��W�����k����1������1�	�t:{�L��S��ǁ���G��*�0؇�"�~&_����<�wA�H|����B��P�z�E~��sB �B}x��73(�R,�fv��(O������ձ�d6�M$�����3�%~��
�vb,ԟ9�Le�)�J��g
�3���˒�S�ca��&:eTW���kÁ ��Nu�͗����Qr��[!���"B�g��{��U!;���?��-�˭X�������U�hMfj�����?��;)\I��A�\UB��F*@f�?��8F^���"�Kb]�n`�)����1Pm�h�SM_�&�֬�1~?��!�"K0p����6����6��[z�;�0дt����JOr��+�|;��-�ޅP��Ʈ���\0���EB-���4A(H�X/P�	�WQx����]'���/��cB���1r�v�p��r~Ԁ"��6���	��Ğ>�9C���#-�'ndN�À�ޯ�u�aW��s)ٯ�.۴�9fA��7^=|�d��[��B�A����Qc�wqq�]���]82L0���� ;�C!�vM�Q�Ԙ�f�i���v5ܫ�����9<�|�q"do�;�����b��FP1�^n�����F�j�!���3�421J���IWSШT���p�IDA��L"o.ZU�C�1�ȭV�j��f�vZs_����W~�m�c��\�y�Fz�U٬��u {@{�ٸ���'�vL.�0�P��+0�(HQ�S2�`���K����0���Fx�`i��e`\��s��92M�V�@k.��I�����s��9X��kH�6l/}* 9Ot%@a
�P+~&u;TYPxQ�Z@H��J@J_^Wא���р�\*�4?�t6��0}-�������|�ـ@��\�%���i��B����UU�l`�����Q�f�����؈q�&R}m�}�����h��HGԲc�mq}�L��+�����b��n=�@ؘ�L �RC:���'��`k*��0C)����:��]@�
��{p5Uz�>��񺯎'�쥴�W%hb���-Y�X��Ҁ����d�՝��}�MWk�?*+��-s�����ĭ^�s{�� ��Prxy	���P��ifo3r
����S��t� �-^J���K�z"&��t=KI�d��'��l4�2��7TEk���T��zp�OU���1��z����HR�kr�W5U*��Ym�>�r�KĻ��!���㥰[�g����j�񛢷�UD�";��v90�I5�%M�Fg�@��P.e�LJ���ϴ/��q�f���x*r`��p���<Y�F�fl����C#Ю.��ۗ1����T(�ɛ�.�l�L����7���t����&�� �ρ�S��cf.~ߕ���m-�f�k[JL��Й���=�f�� �$�K�!�ђ�_qt�ۆ�E��k+%���W�	���(2?�z�
Z2��ƐN֝��[��f�̒���)Z�~)�#/���?jђ�K�N���j9�L���%˻�M\��+�8$�� �קc3&o	��	�j=HX��^�1?p�������&�~�.F3�
Ϭǆ jt5�Vι�~������
W�c�ْ�R�ひ�l� ����.4���h�jh��. 5/n����Gja�����lGg���c���Z�B�3Q� 9���ݯb!�ݬz���'$�� �D�_�n}i��k_%��}�	��$&�~< ��y�Uz���o�@O�?��j̎�,B��;I�u�RW���0�
o�X���k�����iB=@:cg�p����&0���0��OCR+[�A
���`sV�����Ͱ��:Ơ7~�x��k#�#��K��7�ݹ6�2��E��S #��D<��-�6��A�����[$��P�#{"��9������o�����;��'I�V�T���.E*�P*k�p����l�d�t��B�͜�hKCU���2�*}o�b��ʇ|S��!�4'n͉o�$����-��1j�*�]@B�QӷyoX0T�9��9��Wѯ-Uȭ�t�1X���Yj���k0�# ��ҋ��u _�H�Z5W���q����?�	=K��ƻ=.�g X+��!3�U���*��$���f�� �~�/��^�J��8��
��F�!�d���&����ZA�ߝ�(>�|a%��!���%����BP�25&�v��S����A��zm]�;W4�{�^��9�ՖG)�
>��ϓ.��HU��kة u�X�k�sy�u ���<
�#�s�<��쎐GkTXxEn������M��v@.�r@�NZ&����.���i�ɿ�����&{���k��]܆φQܬ�^���@=@#���f3���*Wp�V�ZBڣ�/�wq�a=40�FF��>��Ɣ���A~��0��>��_�F���!� ��$h�o�׽�t�t��<�^�;ڧ�����%�z��6C����ȪK��ƃ�W+�7�=r�w2s��*��i�3X���>��!��G�2����L&oQ���)��8Z!�����;�y�S�y��3��C=�.}���������R:8�Fu$ړ���\E���9�wn_��]��+X�/�1�xy�G*������1��#��g����WA�!U��w%!xV�B]?�eϾB�'LX���HV�q�H�G�('g ��K�7�zd���Ƙ�zŤ����v��0���Kl%���/�R�m�Q䰘���D�?)�0>�D��bXoǈ��N����A_������I��kyv�v�1����\���K�}tI���I��{�V�3��D]�LhÈ���I��#bIYh,��fēZ�[��n��/�2�-vr�ؽ�jۜ�Y�sp�xC��g��XƐd�X�������!72�º����Pe��vu���6ְ��2R,��щ���`�Y Ա	4�h��C Uz�zg�.�S����R=�{���m$��6^h�9�U{Zw�_���/E���|������Af�Y�"�b�O��XGq,��R[�R�e��u������*��h�<�`�3�/\�s���zE5�֚�m�?��R�USL�����F�]A�������3����/�	���I��2�<��Z��J�$_��<���v�Z�������I�G��-^�I���M�8�n��	�rb�Z��u�1U���ȑ������{�.����9-��N|-��P<?�#�B\5�3�ԛ\�����O˿�:��g�2լ檢��?:�'�)������P��&T1:�T�O*�p-&�#<��1.�k�vR�PD��g�h�&
�����S�C)�r��7�xw�]l�:��x}e���3o;O'�ǣ���s'�+�X���P���e�Ŀ�~e�ڊx@m�sk�Y��?+.���N"����Lz���ޝ3���WtJo;?U��� �E�i^��+�2<j��A\���f@��\}6Y��..���� \�@ k��B����j�~��a��j/�	gG�z���iD�f,�QW��� '���Ь���U��M�ON�Խ��5ѽcd%uou9՟���D�N�~�i}����!5�iuB��v3'�Ѳ�i��D���G!��dz\4]���$�|�Y~̉n!�D�f26i�p��4u���D�Uz�x���A�D��ǉ&	�5f񘣮7qy�aNO3��l_�c�z%�I�Y���8�r9IgbUX�P7�����6���E%���$�RX�R,����W/��R&�Ic��;S*ƽ��=]zV����`�q�d�4�T��@��)��~E� D�S�9����=`�`��Z_�K;A��Cc�������M9���r%4�o0M/	� D�*�V����=���Q�Z�Y ����5<����$U&?���-#��Бr�-�89b�2�x���A�{�Y}���*�V�# ��=@�7���sE�*!��nm,R�6���ȡqZ�o٥;?w�զF�hřV��w�P|�0����p�o�A�o/k弫aIA4}dH�Jy����裥�Li$��}�A�~ZIm.5�O5�1$��6�jc�\ҍȪpJ��ed=��f��44A��=p2+:'����#�4�uk�h���*��[�(�������q?uDx�XU$M�w0�JfF�&��d���:�:B���vƐXQL���Qi�Ok��>�eV��
";3���k���2$X	�A]�F%�#+��pN_�{քip �/����}$��7әU/�#2l�T'�W�Y%l�����R{�_�R�N��	nM���$q��(��p����I��;�9�2}2;kA~��e?��`����}`��8�8��5U�\a�� :���ceb�Tق
���f� 9�>���3~�#"��+���ӔF�u��X��uD�Cbx�܀#�J��Q��I���\�]#�	�ٹ��aI���2��5�ӸR
P�2��#e��tu5;._\aZ`�CN��Xa�UC�T�zd=@k�� ��'>��b��ma8�6�ڙ�2R'�"��H���G�QwYP��ʗp�4S�[ܑ���O�{y�H��֪U������pC���L�k�_�1�.�X���9Ϭ��pR8���\�>f]��<0�-�R#h����Qz�� �����?⪦��LwZ�Xt�����H�S��u�T;��0l�b{��	iۓ��&���+,�
jg!t�ǯ.o��/h'`�a�7O��.Gs�l�� 
���b�`䀋P�
or�$B�<���
I��nй��2/<"���2�d�\���йp���Q"T�#��Fl��v�@��
��TM�~���q�h����'X���,H��1��C�n_��9ٰ.jjR�)��P���$�s���8~h����ÈDf�k�����������*�8/ݦ���^OpY�*`�ӭC�
��G�>�W�y5�T]I����������Sf�s �M:����h#ʍ}HXd�̀�M@Ɍ�D?
aY}m�f�}�M�W��-u���Pv�+�\M������-��+��L�Lݧ?K���p��p��N��2�5���D����n_�!#�������f�͹��O�;.k��-�b�g�!�S�?lȪ�;�Q�A*�X�,�,;!�փ�����ZD��$n�YX��H��.��0���~����b����'��@�� �s�h),jŝLÝz��n��K�-<9q�!5ߠ�����M*��u�&XK<�bޘm��I�<�����w�y-��s�'br����re\&���j��x ��rC�|)|�H�*j�(<�h�j�W�(�"a��+!������Cx��m�dɖ��v�+�s�FD��u�۴����-BΑ�,6�O6'C���9�bZ7�q����K�ue]����N�a]�h�<v�(~'�'�0*�Ůe�*6�b�c���CE����8�)T��Z��1ǵ/�(�A�g�Q���󟔾�&��qMliZ��~
�Tп?!�����0K
��;�)+�'"�w[bt񺲨�3�"~w�K��<��55 _aK�K��� di�Ѝ�;��U�ْ���M!�����-�%��\z$�0��腶��AM�4g��m\H*�d����:"��+Ǝ�'����$��~hgPj�������
ڏ�A*��[�GlPG"iB�r�|�[.uE�ծvjC�d����A���"�������	V��%0M�NM�A�M�h��p�u�03a2oZ ���wG����P>�rT���m���'���[_w!��;`"#6���.$������^��t���4�ʮ�X_�����1@^I�E�,�������Ƅ{�jR��J9�p0�C���]V�.�Q
����ь6����<���A_�)����x�T�3�������Se��|����Ϳ��zdV>�ާw�+��1;���û.w򸔢l'B��&�zS��q\�"��R1�G\ة��B4SN�+&--;�M}���aD�1��܆�������24��U�
>D�_
���!���:�n�2`CQ��ۇ�[�ueI�V��Jd�+Jk��0#ܙ�h�7�I��c9'9�����*�R7�SF����B@� �-�\Y]>�O8z��d����^^ݡ��N	���Pd�~�%�>�� %�OF��鷚���6�a��i�7{���-����kX�v���[h�s?� s��s]�b\!�L�Cv(�p����%a�|	��a.�*
�<��G�¦i??Pëh���r τ�ɍ�*_ ��no��v��k07xG�?=�;�u	,�2�v�y�M!m�P]v� ����˞���4�*L/��5�L �w
�la挏N�U�\SJ���[�*�o�[�h�RP��Yu9d��x�P�.`��6K�V��R��e�/U��j:��s�P@s^��ƺL���:V�x;d^�MP̴s�b�����a�=?�&V��$+��۵��f8�΀ޕ*ak�H  �@&�0��E�(���X��.Y�B=����f �2�AL��	||��"������~���9@˲�̻��d޿l嗑,�	eT�]a�y6|����A1q�Z���JL��L��_բ><�o���
5?�K,�^(��ӥ0�Ѫ�zP���_9���M�n�܉ʧZ�ʯڛ�1Y#��D=P0�����TZ����ZHV�#Ɉ_}��n�m͙[9��L�wQ{K�S7���ʒ�Ұ !��&��0:P���摇3&S�z(m�KW��C���2�Y
Z�8�ټud� �R��磉r�W����~�';A'@{��ϜX�\��HB� �fc뎅.������%J���0q� Ü��J�O.x���_7�i�V��gH�5��7��9G��4�
6�?�sU+w	���ȷ�B�e&�rk�3$V�x �pK��t������W a��|�瘕��h��Z��L[����+��5̖��W^P�����xe3p/k���4a!�gc�6�����������d�P�O5�í;��Ub�ø"P����IC�4GF�)t��A�is���`#%���~-�������TB6ְM��,w�h�|���`�U�X{>�Mؽ�f��^$@>�e_����Ͼ�®xM��/�.)�{w��a4-;���ӦoJ@�0�í���{�]�X��\Ѓ���Wn�uz��,RƐ0��ՔqdtkgDX4��Q����O�����K�<RK�rb0Gz��|���={/���,�N�QZ��Q�P7�#��|�>���WW8�E��q�։���r4?�xITG�.�>�ݙ�S+[�T���ͨ�Ȏ��]�t��͇�7���K^J���F�1d��Zx*9d��LՊ˩~��0��w�����j�q>����(?�TQU�7�AK,)J��6��8
C&��5F;��뽺��T�I���6SQX�������%8�:An���k����X޳��ҁ��R\�~MB�3�7��hg���(�i3���k` 
:�xgmq�s)��ĵ��f�S��Y���*ҳU�Q1�C��V�/���\� )���d�m�s.,{�6��8g�M���/zUE�$̦<�5��X��:�����H���*'�yEM��qG�[E�pN�Fv*ڣ����9�������Α�/C}%_�gMGB�l�XuW�h1�qN�ꆭ�e������m`r�Ji8�@������7�V����s�W����b��$�B�RE*_��-����t�a��hDA�6E'�I!{|�Q�r2qaC��;8U�$�:�-��Ddo�A���@@�?�K���s3��K��apW����<�u�&��̎�����<2���s�����@o��q�Y�V�f%ߍ/<MK�9�4�)	�j�:��-�>�B^<��pѵ��G!�C�eş� �ُ���d+�>�H3	H(�[��FM/��(4���"�!Oʴ�����p�u)�83��6��(�C"c��MuY�.���74W�m�,d�����{��\韮��~Z~�0�j�>a}�3?~1+V�/Jۙ�y�lծ�Q�3$Z @N%�C6�e�3�;�+`���I;>��! ��O9{��L����J��+�?2&*��*Ƚ�C���R�rd�C���N����� �拯�����ILx�)h4��� [N��V���M�L��(��nL���FO[�#���� b�\�J�&�Z��|9��1C�=ŀF󣂀uY)$��D:��Q�7��˕�T�%˪����<Z�RcS��r��]�NycЂ�!�4��s��^�BNyDҎ��d�Ӎ�M��Wa`Xb}������\�.�������vn�sDq���z@�u�`��zӰl�޿���:¨5��xmL�v-S'VZ�^�Z���6���i,Y�� 0�$U���.�);��Y��Wq��t���]���E��B���JD#��?��fd���D)�4�*����49.-���c�l�![�w�?o)��1fv;�P���'����\5B�e�q{�9sĔ���S)�M�Իu�FYr�A�T��h�q�N����1�*`��v���?HcHc��$w�h���l�4lqSx#�����'rw�t�JFO����V\�|#uޡ��9�f�V~���w3|�3�L�_"�19	�����d?��Y�$�������gi���*��c������CF�7��I�)PZ���x+Β��[��85�.%���B<��6:Ѥ i-i*���oL��.��vp6�~���Jg�W�H�l�|a+�Σ�	�"1�̡�-(��&��j櫸p�`d�>��O%ν0NT�'/be��	������ο�\�J�ë�����?Z���1A0ED�Hѥ:��N���|�^X�8l��Y"&
�0#2-��G6peAF-��1�Zx�r��з�{��h\{i��rK�>�/�A���3�Gb��G��'s�n��Iz=�B�����C0�����xp��S��wԑ�}~��i��T>I�!�y���΂��8���.V��V��O���`�<k�xJ�T`颧����=�d@^/�w{0?/�یӠF�tg)y��[�9��2�����,P���\��y/�4!h�8y���*����.���/eشC]1F� �w�a~����ic󔿽V�\�7j�K�I�&��x�@$Q�w�Hl6���dk#�C ����`�(�y�o�i5�t��.�GhU�x�O�|��X� 2���v�������&�K���>�RN�Tc*�P��RjF��V�[��r��¿]���HйN-tN���V;�G��^<���_��S}krq�"X{?|0'>�5�u�u���A�q�P�,E�{�d�%����.��1�2W�t�c�A#�sn�gp�gR�v�څ-(q�W��ƛ�����8�.�9�6� e����g�p���T]�
/%�c`Q���'z��=���b��뫃��/�5�:5�O�mM�B�u[.���ܥd<� ��y�8Z1h7w�5�?��yeFt^�콇ݸi�L~���f 5��A�@0���C������//}��V!D}�'b[|��hnN�X�t3�+��@��	�X�65g�-����#4 6��N��g������Glf0������Rc��LTx���Yߕx�|_�j �M�(�1��±9��:q�ŧ��?��;����K����Y�
��o��f��}Z����^L�?&�y�z��|��7�р�'�x}Yb�X.մj����l���wzj�n/�2��蹠���RZg�tG�8��%yR�%��i>�C��<�HF˝@�0�m�ᥖ`��pD3~r�K�g���,C	T�h7������O"\q��m�$���~�җ([������<ȯ�$�T�bl���
�����N�sx�]֕:�G�E3^Rz�n�$��?�F80���ط$��d�D;K$*2�sI��Q���~�Y�(J\��j������	���j������0��X��k���5+�����Ed'�&"X��?&sSy�8� �̀�2��gL���LN"r⌮6����x��`w*���3W7fC+���=��s��}}]"G�d<�$Dw(W��y�I ����]`�g5��7I��WR���t���Sxd��d%���,�v�P��t��O�+��xQn!�B�z;O�۸P?�b<:fe��������d�s)''�/�����d�XҺ�Q�J���6��si^�U?VڈU���;Hޜf�� �'ˣSĚd��ܴ��H8�l#:_J�8��Z�q��j�n��
C�7�	BT���w����pi	@͛+�Z�[ʀ�t���(�hTX�P�W���a��Bَ����l_F�.[�,�h���Z,�uo��Y5-ns�i�igxS��8�*H �%��fL� ���/�;�%N,\����O�j��r�uV�4�����T��ض=ߕ����
j�A�S%�X���	��l��b���~���-������K���C�fr9~ Z:I�9[.�8�N`�&�gH�fL���顫�7�uԄ�{86�q|):i#�//��L��&�'@��v�:�?�-L��+ɽ��yE�VdY���Y�{�Ä�'-GXB���n��D㋚m�3C8�����ʒ���3��Ι�}4!u
��xħt2����{d�-�!�eM_���W��8cP�Rs�����M.�;�@�4&��� d�@/ZC]��Х���q�ЊxSp 9 �MP����}� �2*�
�TI�Yœ�����6)9��s�0~eS��aj걍�-ھ�b��D�K=�:�ݝ%��paw �����ׄ�S��&�'��*�W���.�78��'�a�k��sf�B���@�PE)£�\���Qb�"��k��97D�i��&����<���z��=�A�6��W���"�Z�i�֟��.��;j�no��Rl�p�ڗ�;�G{{���/��c��)M%�\ h,UԀ8=�DĹ�Қ8x�LL��y�,����B��<"R_1�5����ۑ��M�B��j��(xA�s�J�Z���A��y"��nE�f���Й[)K� ��|^�Y�ѪW����,�w�n��ӗ(�	�d!�����I�/e�LE��S|���ĥ���zL�� ��,��������a���K�E�����n�T����d1��.VLA��OE�	���J��B�a���\�}�+ݒ8�ոj�c�,�N@��e��0�KזϚ���!㚥j\��YaJn�Bh'%�p=�n	��	�d$L05᭳�_!� �9�
�h�oPB[t��r�ϫ|�u8��8�����`���#����x�<�rX,�X��������VK�t��GdQ%��^k�X���P}m���V�*#���zJ	$�y�B���躉�g���8�v��k�:������n��f�LK�������qmGC�,W�p:�j����ŨV��� ���Z�J��
G>��;7��nj �Z�(-4o3�g��;�����!�<���yTT
[���=��^@�����x��ǽ�w�L����s��ķ��*�Ci(�9�K�^�ѯs�ĺ�h�0�^�[�Ō$�Xf��d��!b�1}���X��׉��4����&R-�V�4ո�E�x���#Ɲp	��x���_!���+�Ïk)`V#�/������@��X�<
�XX[�2�e�	���(���i�Nh2_}�k ,p���^=�j?m���h+p��� F�V��p�P�X�AN��*�Cm�H���rkNe��y#�ǆ�+ߍd�V��㚀q�J�H��� ����`6�j����y���$r%toD(~H{]
iPs���,q��}&�xmN���V��xAS�,pa�Bj�{�"��2���l�[ �zr3���B����z2RIO���'|Jc
���#a�	\0	��kѕ��|g
��Z"9?r.O��]��=�l�i{c!��=Z�x��
{�7���B���������Sd~�z�p���i��״�����a��_k��c�b�6p�i�)�9��]���?�l(��A]�wr�������X�*�瘌"�N���(�v�"����/ҸK����$/}ިd*�P�{�A ��w�: ���NQ��r�,v��Y��U����V>�5�1m^����'�⦇���I��
@mC��a�t�"���qSk��x��R�d7�T�(9��ߕF�k�d��3�K�O����l�֫��Hu��X�@��t:,?��0��v�6�WG���r��-����&8�;���޳7�H�!�����{{����5J���#HC��5@�9Z��]%���'�G5�%�I��\i�����D) 9B8~Qq�S��FiH���T�r��A��Ut��E���{����¤��Ť���!o\:}��əN5���:̚�_�m���q�B܃�EN��;�o$.j�{1�U�#vS��r"9�����;�l��&�f:�)?ez�)�\4G���ݿI�I}6�Xn/�=l�	���d���v�|t�AY����ω�	2$��豔<BA��O~�&v��S�2�`b�9�[�bp/�	k/�d�tpg�/�^E�Z:.���/7H�Yu�D������>t�����O~� 73�����U��I��
͓�^7��=�̗b�!}� �{�����?fJp�*���Ƒ�B��ouɶ�p_���"��}a�~9#wwA1��pE��bL3��W�5�pXJ}6A����K��*>�6S��Sۘ�w&��W��4�|8ל�x�U��{1B�Pdl��)�y|��k��ٍ,��f4#4�g�tάK�LEp[ B���=<��Y���a��hi;A�5�.��[�A�`�)�]=�9/�5җl���>�fȭ9�9�%_�}��۩��f��J���[�(�\�
���Y�ѳ��{��)WQ�^Ⴕ��Q�R@���}�[�i��$-L��������+��m��t�X�*`��_J��4ıw�|&��/e������-#Y�9��G���'���V���;z�hU�PR�Z�9�o�w��>���ϊ���������	;e�`�����D�\�7U�q6
���0D&�Z�H롡w��X�|J��%�l�Z_:�_n�?��|�����1Z�G&�])�R��g���`�yt.�Ry�Pa�j�n�D1%�19^g����u��1ꃎ�ư���o�a��kUs��� �)L1���i�D,�ړ�l����K+-sP�Ew�[����{<����������g�d��΢�;l$i�hc��-�>k������'ymyOk��A6��{	��g��Æ@�z�`���b[Z��M��喝�Z�.]Fr���vvA�J���iJ��~Aaן�R��\ނ*!:�N�ɳ�.��a�k�\��n86�+ S�(��(D����dlez��֡h�J��E� �v3���s�S^^ړ��OѤCˇ��Hг�wg�
���Ԉ�nS���뾋���R���tS��&t���a��G���-�Ak�n&?1[q�û#{��s�a8�ԫ�K]Y������� 4�~�6m��w�!������mm*�ǎ��^��۷�t?��U��бv�7o4� ^k4�P]�L���U�:V����r麹�9Y���10�J��Ipܙ�'�bzqt��g-
�l/=Ѐn�����ѳp'�O�1B$���d_�'�pI��g��؈Y�
�>�Vw�"F� 1)����=�ڂ���I��'e��`�o�?��f�\_�Faӌ�:ڔ�4��iVB\��`���݁'�raP_�_�XT�[
���mBK78{�'lAbu<퍨�S�o���/ ����6����(*��qbJ8;��~Рu?a�8� ������ɔl��j����O��Et)RN��s�c��&p5h5���}��1,�\��X���בf:���|��8
�1�����{�\� Ѿ���G�69���m\��e�N�y�$m�w4+�����3�\�,ՄIbT�L �|A~N���~����A����ĕ�}~}�f�A���iU�2:6�d��8��J-)����ժ?��.0p��A��&>�a���Őf=-}�얾�oh"6뺾xa~�V,ٻ��O���oHܒT�0 ���P""�;Y0��w)(�P@r(�m��"<�LE[7��_uU��Ҧ(���I�T|�Em��@�5`���_��=�_
����g�V����C�8��V�z[�׍�5j��)�p�^M'�֝��f ��1������RY������%�@}F���`��h����V/>,��$���zB�b���\TT�9>�i�%O����\:���e����/��I*�W��ScX�V����%�籖����ғ:)	�ay�i���	YON9NVi��Y�2x2v,%�g�̕����=�Z�N��QI��_�(�������{�%;'��\	� /2>�=e�q˖�h��E��^J�툊Iߡy ���;6�d�Iw,�X��t�4�<3��b)�r�C�՝� $�[�eP��>�g�2��5x�Ǌ�.F&Ԫ��'M�FO[��z����/dB����.x�~ ���w^����<َ�志�`�Qi�Y�71t�8H?ޗ��`�"'�EX̥��t�տ	�ha&cq)h8�v�\���P1"� A�����]���3٫��~� N�n8��{�6�=����nZ%����g(�P�MK\v� H]�>@��B9�ԟ��'!�ݒ2��ly��}�|��pZ4��%����ӹđ�>���v=ؼ��p�]���a¤z��x�7>�?}$6��6�z�a-���ʍhϞݏ�����\I'�:^�^6��]#E�!f椒��p[���I��