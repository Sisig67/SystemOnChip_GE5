��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�H�u�%XPcr{r�mO���2i��'�d�A�I~[�"�մڎw�dj�o�v{'���K)s�솱���4W��%�":K����;�;�Y�g�?��X�af��H^�c^�)�Mz7��֜$+�0�\���p��R��0��3���O5����+LB�¹�+�X ��`4ɞr��<:�'�j�I��<�[�;6+JT��/��z��Z�b��jBuP���(�w���ət�'�<�(_�l��)s�R%�%�R��о�ׯO;�����k���!Z��^��B�x%a:�b�Q_�n/�*��"���^[�e�3���UZ(`S�st������'�@�Z�f�UAL`Y�7� �a�j���'���
�4�!\r������E��0.ۢ���o��:�k���:��v��kU;*��(zȩ�Һ8��Lt߶Ţ��{�~5���c8z10 &��\"/Rl����R݂r�d�m��)�*�/9�_�S�P���e��1i{��pN%�� �h���6���%�ڃ���Ƥ/0������n�2�km�	���Þ�����<g`>X7��Ǔ��B�@��pu�������$�#�]��3QX���/h��k�Ź,S6ݓbyn/�>���x-���@%qs5^₽�Ą�|�EKt�/���������Pd�L��Tb�Wz|R�ך|�T_����ٜ(���s��쥣'�s3�u��|n���ӗF<.���U��D��f�r�u���!���D�E�S���0'��C�[�#����Fɡ����%QN������/����a���G౰�!�_77��HC��x����\a��\>�J��l�|�c�ME+�x����}�H�;�2VfjmH��0u���ԝ�O�z�G�P��{�H]YVs��e�,���|�;e.�,_W��J�L�:���My��E��t-'���|��%�W�Nus2�r�VNy�t)`������p� ^�X4�nh	h�!}J��'Fc��$`yµ_���5W���L������^�Xz���:QeY�sU��\6{wA�^o �R�D'Y��ZY�J�'�BYKF������� A6�vH�P�t�!4�ʨS��ɟ3i����% 8��U�T�( ��?Y�_���u t��ߧ�B�� ���b���$�u2���Z[g+^;�c��|LJ�ٺK�s�'����8?&m7���هV3Uxe�C���~��4�K�2�=�����D���{0���"g�R�v�9~Į����07@�p�S�C��.	
�
��ӫ����A �)�me>����LU��g/�	)c?�~BD)!;����s��U�c��0����<�x���@�$��lT������Ѱݷ&a�Qc�M��U�J��Sl�9��~���ZGG�q�0�{;w���O��
���+��T���N?�Vo*l���
y��P�*�L�\�pY"J���0Z���|�ٟUӨ��b�����e�!�g�J��&�9Ki������J��ƒޜ���G�E_���5�0��觲�3�#.#\  ��ܢ��H���N#Pm����tz?e���Y��Vw�+ "�+ڛ���>R?f�M��&A��������(g��_���p��%L�y"�h�2�p���K<�[�؟m��������L.dܝ�҈Ѻ�G���/f�^���»�ڕs�f��zT8���1$%F?IX�{��Ͱ:i�F�7p��RN?ő���
�ὼe�$Xi�(�)Z�ſq"��R��Cl�ߦ�7��Ё�Q�>�%�5��� ?�˱^�V��!�_�SS�|�*��%a*�y�> �	�;��F%gc�̆��1�b�_2ϼ"�[`m��7���1��=�3�>z����˨!J#[��2�GY��4��vJ��誥У��KV��Q��_�I��Zb�F��4�SU�>�|��"�F��F�$�j��ԗS8i>U�![���
u�]��#�&ٶ���F+�e`5ڭ���**D��&�k�鐿Q��R�ܤ"(�
*�}.H�^�����6(:��s.��e�G]U����	��d��Ӽ+��^τ��*�ҹ���Lo��d��L�� �$t!c|�f=r�:��~ՙ�1 }�(%�]BW��%ԡ��:cK6ҍ7;��1$ٔ�@9e��랶N����_؜CW}~2y2�Qp*4��3�G�3��	r@O��<0'�F^Q��xe��~����v��׽;��P����+�+UEV�7^����@��}~�]�����_A!fv]dTCN`T��̎��-�M[K)BmI`π��7�����(Ӌ���4��}��M��uo~�l��\WW$��(Q��f�^���-�W0�'�s^1�1�rV٢�/P�G
���������w����Ϸ(a�4�&}�"��[P�C����&ֈ2\#J;�Xf�R	*��uc�>?�{��ID�G�'�ܶ���{ _�d�/6��q��� ��3#�'�ߐ5�wvz����H����}�oH��X��έI$�IJU�d{�CT~F�G*����$�R1P]��":/S�^����T�ӈ�'	��{�7v���;,���A Q10n}8D��I�2�`�a���������e��G�_hA�$�|�(���A��1�w��'��'�Uy\�5.h$���D��h�Ԇ��_��(�āɦ�Rp���%[IE�Ou6)Ws�GY?�R�BȘ̼P��	7�S2�ꨅ/���H|���ho:tcX+M�U]t�1���M���yt�x�j��6mv�v=(�����72`t7�츬Yab�C�(�qdR3�1�0#!�N
˯�8Pl;���`s�b�$�j�i�	Q�c���ed�ʝ�m���4TT�
�fNte�m,k9��'Y���&	�Nz5x*�N�)na���حl�U��v��9ut��u���ӹ�B��$�Ј�LD���qp�K�F$�������R�UqB�}�֞L�_�Tю	KX�`N�pp��Mߊ�F�|6����&ld�=1��x�%9,�m�'3!�L��
��Sdt3���渊�<*ԉB�V:x�|��������㪬;xN�v���Z�gaѢ�"�1r3�e�9��\�Ւ'bpP֪G�ɑ�
�r'���k���zX��%�I�qM+5����D�⑑��.�<���*�<�0:h�u��ޘw3��$8�!����@N
V ^Q3�(���x�9���y`����ARն~��v��P��W��v9��I��� ���y�ܧ{4iLM���9`�{?*&�����d�+�T'��%Ck���)������l�}��3V �S�֝$G6l�"g_X��?�/g�߀Vud9E�mR�.�+��������Ӌ���eQ�t��R�J�����}�"��,(�)Di��m�S��ݨD�R"2����D�(��&�� Jl �h��5�T�>���Ok-�
y��\�p. q�u4J���щ1��bCU�n�e��_U�ɹH�s������t��,dB��_)�q��~X�Zʣ!:@^�G]�WT��4H�y՜��)���6���b��.�� ���VBL�%l�㌷a�������6*��;��b�N�{��5 �Vu����2g�V�	&�>'�~�9�p
q��G���f��z�/3�oQ�}��t��5)��D������(�-�Nld��d�Y��v*#��D�5��Tc����u��p�	��A��z[��u�����ޯ��E���^ى�	vx�T7$�ٿ�Ն�r];v�R��-�2�ő'�[j�@{� �/��3j�����P��N_'R[0�de�P!�*�̋�-"ʭ*逊����6N'_M�8�L��P6�n�mG��c0 �����u2H�L]sė�u*����� S�N�t(�T�8�^�w�8��v��>|��p��Ȁ�R23�M|N��ݵ�ݵ�ӷC��GZ6���i�9L��y��Dc�h�#�w��p¬�1�a�?2�D���f(�l2=X�<�!�W�Ps @���mX�ł�K���6����.u���y�ܛ$��ȋ�����O��7Oӄ����Bp+ܷ��;�i����:�uƋP��+ "@����Ap�_&vkxG/�(����bonI���+��E��۴XTJw�.i���΅?	���WʒIB���RA��y�R�򐣎�k�Z�j�pA�H9��5�}yeڅ����WZ��}*��f;�,�Ft��j�`����_(���9�ez�>����egf�K����sn����>-�j��i5�r��ҀC��ĸG�}:$������Wf��玮J��7#�Hqh��Ź����^�%�§@�!4�����
�j������P{H-8�5�#�n��S�6:��y��/mL�x����5��%a�;��;"ZJ��G���k�灑n�p�nC���'49:�p��Ҭu�b`t3hxԧ<��:r{�#�-�A��b�Q��>@n�U��쾚��kx�U� -�3/Pg����s��� ,���9�_���5Y�d�#޵!�gy��E�� ����x�U���TxIn�p��d�0�U����C���"MĀ�'��!���j��Uj	�����v[e;�xpb�/���Hu�E@�N�o�6�L�VQ� Қ��-��륋ݹ$��A��e�i